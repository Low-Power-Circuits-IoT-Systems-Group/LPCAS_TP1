magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< nwell >>
rect -201 -36 119 236
<< pmos >>
rect 0 0 30 200
<< pdiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 151 83 200
rect 30 117 41 151
rect 75 117 83 151
rect 30 83 83 117
rect 30 49 41 83
rect 75 49 83 83
rect 30 0 83 49
<< pdiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
rect 41 117 75 151
rect 41 49 75 83
<< nsubdiff >>
rect -165 151 -107 200
rect -165 117 -153 151
rect -119 117 -107 151
rect -165 83 -107 117
rect -165 49 -153 83
rect -119 49 -107 83
rect -165 0 -107 49
<< nsubdiffcont >>
rect -153 117 -119 151
rect -153 49 -119 83
<< poly >>
rect -18 282 48 292
rect -18 248 -2 282
rect 32 248 48 282
rect -18 238 48 248
rect 0 200 30 238
rect 0 -30 30 0
<< polycont >>
rect -2 248 32 282
<< locali >>
rect -18 282 48 288
rect -18 248 -2 282
rect 32 248 48 282
rect -18 242 48 248
rect -163 153 -109 200
rect -163 117 -153 153
rect -119 117 -109 153
rect -163 83 -109 117
rect -163 47 -153 83
rect -119 47 -109 83
rect -163 0 -109 47
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
<< viali >>
rect -2 248 32 282
rect -153 151 -119 153
rect -153 119 -119 151
rect -153 49 -119 81
rect -153 47 -119 49
<< metal1 >>
rect -18 282 48 292
rect -18 248 -2 282
rect 32 248 48 282
rect -18 238 48 248
rect -163 153 -109 200
rect -163 119 -153 153
rect -119 119 -109 153
rect -163 81 -109 119
rect -163 47 -153 81
rect -119 47 -109 81
rect -163 0 -109 47
<< end >>
