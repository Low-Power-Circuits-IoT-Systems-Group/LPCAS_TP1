magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -17 -17 17 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -23 17 23 51
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -51 23 -17
<< end >>
