magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -17 -23 17 11
<< viali >>
rect -17 -23 17 11
<< metal1 >>
rect -37 11 37 17
rect -37 -23 -17 11
rect 17 -23 37 11
rect -37 -29 37 -23
<< end >>
