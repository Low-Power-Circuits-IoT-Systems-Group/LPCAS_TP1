magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -45 1329 -37 1363
rect -45 1261 -37 1295
rect -45 1193 -37 1227
rect -45 1125 -37 1159
rect -45 1057 -37 1091
rect -45 989 -37 1023
rect -45 921 -37 955
rect -45 853 -37 887
rect -45 785 -37 819
rect -45 717 -37 751
rect -45 649 -37 683
rect -45 581 -37 615
rect -45 513 -37 547
rect -45 445 -37 479
rect -45 377 -37 411
rect -45 309 -37 343
rect -45 241 -37 275
rect -45 173 -37 207
rect -45 105 -37 139
rect -45 37 -37 71
rect 311 0 330 1400
<< pwell >>
rect -71 -26 337 1554
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -45 1363 0 1400
rect -11 1329 0 1363
rect -45 1295 0 1329
rect -11 1261 0 1295
rect -45 1227 0 1261
rect -11 1193 0 1227
rect -45 1159 0 1193
rect -11 1125 0 1159
rect -45 1091 0 1125
rect -11 1057 0 1091
rect -45 1023 0 1057
rect -11 989 0 1023
rect -45 955 0 989
rect -11 921 0 955
rect -45 887 0 921
rect -11 853 0 887
rect -45 819 0 853
rect -11 785 0 819
rect -45 751 0 785
rect -11 717 0 751
rect -45 683 0 717
rect -11 649 0 683
rect -45 615 0 649
rect -11 581 0 615
rect -45 547 0 581
rect -11 513 0 547
rect -45 479 0 513
rect -11 445 0 479
rect -45 411 0 445
rect -11 377 0 411
rect -45 343 0 377
rect -11 309 0 343
rect -45 275 0 309
rect -11 241 0 275
rect -45 207 0 241
rect -11 173 0 207
rect -45 139 0 173
rect -11 105 0 139
rect -45 71 0 105
rect -11 37 0 71
rect -45 0 0 37
rect 300 0 311 1400
<< ndiffc >>
rect -45 1329 -11 1363
rect -45 1261 -11 1295
rect -45 1193 -11 1227
rect -45 1125 -11 1159
rect -45 1057 -11 1091
rect -45 989 -11 1023
rect -45 921 -11 955
rect -45 853 -11 887
rect -45 785 -11 819
rect -45 717 -11 751
rect -45 649 -11 683
rect -45 581 -11 615
rect -45 513 -11 547
rect -45 445 -11 479
rect -45 377 -11 411
rect -45 309 -11 343
rect -45 241 -11 275
rect -45 173 -11 207
rect -45 105 -11 139
rect -45 37 -11 71
<< psubdiff >>
rect -45 1516 311 1528
rect -45 1482 14 1516
rect 48 1482 82 1516
rect 116 1482 150 1516
rect 184 1482 218 1516
rect 252 1482 311 1516
rect -45 1470 311 1482
<< psubdiffcont >>
rect 14 1482 48 1516
rect 82 1482 116 1516
rect 150 1482 184 1516
rect 218 1482 252 1516
<< poly >>
rect 0 1400 300 1430
rect 0 -48 300 0
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< polycont >>
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< locali >>
rect -43 1516 309 1526
rect -43 1482 8 1516
rect 48 1482 80 1516
rect 116 1482 150 1516
rect 186 1482 218 1516
rect 258 1482 309 1516
rect -43 1472 309 1482
rect -45 1363 -11 1400
rect -45 1295 -11 1329
rect -45 1227 -11 1261
rect -45 1159 -11 1193
rect -45 1091 -11 1125
rect -45 1023 -11 1057
rect -45 955 -11 989
rect -45 887 -11 921
rect -45 819 -11 853
rect -45 751 -11 785
rect -45 683 -11 717
rect -45 615 -11 649
rect -45 547 -11 581
rect -45 479 -11 513
rect -45 411 -11 445
rect -45 343 -11 377
rect -45 275 -11 309
rect -45 207 -11 241
rect -45 139 -11 173
rect -45 71 -11 105
rect -45 0 -11 37
rect 0 -48 300 -42
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -88 300 -82
<< viali >>
rect 8 1482 14 1516
rect 14 1482 42 1516
rect 80 1482 82 1516
rect 82 1482 114 1516
rect 152 1482 184 1516
rect 184 1482 186 1516
rect 224 1482 252 1516
rect 252 1482 258 1516
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< metal1 >>
rect -43 1516 309 1526
rect -43 1482 8 1516
rect 42 1482 80 1516
rect 114 1482 152 1516
rect 186 1482 224 1516
rect 258 1482 309 1516
rect -43 1472 309 1482
rect 0 -48 300 -38
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< end >>
