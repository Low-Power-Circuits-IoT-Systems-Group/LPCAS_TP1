magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 600
<< nwell >>
rect -47 -36 401 636
<< pmos >>
rect 0 0 200 600
<< pdiff >>
rect -11 0 0 600
rect 200 555 253 600
rect 200 521 211 555
rect 245 521 253 555
rect 200 487 253 521
rect 200 453 211 487
rect 245 453 253 487
rect 200 419 253 453
rect 200 385 211 419
rect 245 385 253 419
rect 200 351 253 385
rect 200 317 211 351
rect 245 317 253 351
rect 200 283 253 317
rect 200 249 211 283
rect 245 249 253 283
rect 200 215 253 249
rect 200 181 211 215
rect 245 181 253 215
rect 200 147 253 181
rect 200 113 211 147
rect 245 113 253 147
rect 200 79 253 113
rect 200 45 211 79
rect 245 45 253 79
rect 200 0 253 45
<< pdiffc >>
rect 211 521 245 555
rect 211 453 245 487
rect 211 385 245 419
rect 211 317 245 351
rect 211 249 245 283
rect 211 181 245 215
rect 211 113 245 147
rect 211 45 245 79
<< nsubdiff >>
rect 307 555 365 600
rect 307 521 319 555
rect 353 521 365 555
rect 307 487 365 521
rect 307 453 319 487
rect 353 453 365 487
rect 307 419 365 453
rect 307 385 319 419
rect 353 385 365 419
rect 307 351 365 385
rect 307 317 319 351
rect 353 317 365 351
rect 307 283 365 317
rect 307 249 319 283
rect 353 249 365 283
rect 307 215 365 249
rect 307 181 319 215
rect 353 181 365 215
rect 307 147 365 181
rect 307 113 319 147
rect 353 113 365 147
rect 307 79 365 113
rect 307 45 319 79
rect 353 45 365 79
rect 307 0 365 45
<< nsubdiffcont >>
rect 319 521 353 555
rect 319 453 353 487
rect 319 385 353 419
rect 319 317 353 351
rect 319 249 353 283
rect 319 181 353 215
rect 319 113 353 147
rect 319 45 353 79
<< poly >>
rect 0 682 200 692
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 600 200 648
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 648 50 682
rect 150 648 184 682
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect 0 682 200 688
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 642 200 648
rect 211 555 245 600
rect 211 487 245 521
rect 211 419 245 453
rect 211 351 245 385
rect 211 283 245 317
rect 211 215 245 249
rect 211 147 245 181
rect 211 79 245 113
rect 211 0 245 45
rect 309 569 363 600
rect 309 521 319 569
rect 353 521 363 569
rect 309 497 363 521
rect 309 453 319 497
rect 353 453 363 497
rect 309 425 363 453
rect 309 385 319 425
rect 353 385 363 425
rect 309 353 363 385
rect 309 317 319 353
rect 353 317 363 353
rect 309 283 363 317
rect 309 247 319 283
rect 353 247 363 283
rect 309 215 363 247
rect 309 175 319 215
rect 353 175 363 215
rect 309 147 363 175
rect 309 103 319 147
rect 353 103 363 147
rect 309 79 363 103
rect 309 31 319 79
rect 353 31 363 79
rect 309 0 363 31
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect 16 648 50 682
rect 150 648 184 682
rect 319 555 353 569
rect 319 535 353 555
rect 319 487 353 497
rect 319 463 353 487
rect 319 419 353 425
rect 319 391 353 419
rect 319 351 353 353
rect 319 319 353 351
rect 319 249 353 281
rect 319 247 353 249
rect 319 181 353 209
rect 319 175 353 181
rect 319 113 353 137
rect 319 103 353 113
rect 319 45 353 65
rect 319 31 353 45
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect 0 682 200 692
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 638 200 648
rect 309 569 363 600
rect 309 535 319 569
rect 353 535 363 569
rect 309 497 363 535
rect 309 463 319 497
rect 353 463 363 497
rect 309 425 363 463
rect 309 391 319 425
rect 353 391 363 425
rect 309 353 363 391
rect 309 319 319 353
rect 353 319 363 353
rect 309 281 363 319
rect 309 247 319 281
rect 353 247 363 281
rect 309 209 363 247
rect 309 175 319 209
rect 353 175 363 209
rect 309 137 363 175
rect 309 103 319 137
rect 353 103 363 137
rect 309 65 363 103
rect 309 31 319 65
rect 353 31 363 65
rect 309 0 363 31
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
