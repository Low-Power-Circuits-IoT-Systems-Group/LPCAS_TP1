magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -160 26 160 27
rect -160 -26 -154 26
rect -102 -26 -90 26
rect -38 -26 -26 26
rect 26 -26 38 26
rect 90 -26 102 26
rect 154 -26 160 26
rect -160 -27 160 -26
<< via1 >>
rect -154 -26 -102 26
rect -90 -26 -38 26
rect -26 -26 26 26
rect 38 -26 90 26
rect 102 -26 154 26
<< metal2 >>
rect -160 26 160 27
rect -160 -26 -154 26
rect -102 -26 -90 26
rect -38 -26 -26 26
rect 26 -26 38 26
rect 90 -26 102 26
rect 154 -26 160 26
rect -160 -27 160 -26
<< end >>
