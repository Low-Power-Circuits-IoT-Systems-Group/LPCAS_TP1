magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -26 26 26 37
rect -26 -37 26 -26
<< via1 >>
rect -26 -26 26 26
<< metal2 >>
rect -32 -26 -26 26
rect 26 -26 32 26
<< end >>
