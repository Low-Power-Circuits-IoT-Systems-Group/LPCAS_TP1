magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 0 0 19 1400
rect 337 1329 345 1363
rect 337 1261 345 1295
rect 337 1193 345 1227
rect 337 1125 345 1159
rect 337 1057 345 1091
rect 337 989 345 1023
rect 337 921 345 955
rect 337 853 345 887
rect 337 785 345 819
rect 337 717 345 751
rect 337 649 345 683
rect 337 581 345 615
rect 337 513 345 547
rect 337 445 345 479
rect 337 377 345 411
rect 337 309 345 343
rect 337 241 345 275
rect 337 173 345 207
rect 337 105 345 139
rect 337 37 345 71
<< pwell >>
rect -37 -26 371 1554
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -11 0 0 1400
rect 300 1363 345 1400
rect 300 1329 311 1363
rect 300 1295 345 1329
rect 300 1261 311 1295
rect 300 1227 345 1261
rect 300 1193 311 1227
rect 300 1159 345 1193
rect 300 1125 311 1159
rect 300 1091 345 1125
rect 300 1057 311 1091
rect 300 1023 345 1057
rect 300 989 311 1023
rect 300 955 345 989
rect 300 921 311 955
rect 300 887 345 921
rect 300 853 311 887
rect 300 819 345 853
rect 300 785 311 819
rect 300 751 345 785
rect 300 717 311 751
rect 300 683 345 717
rect 300 649 311 683
rect 300 615 345 649
rect 300 581 311 615
rect 300 547 345 581
rect 300 513 311 547
rect 300 479 345 513
rect 300 445 311 479
rect 300 411 345 445
rect 300 377 311 411
rect 300 343 345 377
rect 300 309 311 343
rect 300 275 345 309
rect 300 241 311 275
rect 300 207 345 241
rect 300 173 311 207
rect 300 139 345 173
rect 300 105 311 139
rect 300 71 345 105
rect 300 37 311 71
rect 300 0 345 37
<< ndiffc >>
rect 311 1329 345 1363
rect 311 1261 345 1295
rect 311 1193 345 1227
rect 311 1125 345 1159
rect 311 1057 345 1091
rect 311 989 345 1023
rect 311 921 345 955
rect 311 853 345 887
rect 311 785 345 819
rect 311 717 345 751
rect 311 649 345 683
rect 311 581 345 615
rect 311 513 345 547
rect 311 445 345 479
rect 311 377 345 411
rect 311 309 345 343
rect 311 241 345 275
rect 311 173 345 207
rect 311 105 345 139
rect 311 37 345 71
<< psubdiff >>
rect -11 1516 345 1528
rect -11 1482 48 1516
rect 82 1482 116 1516
rect 150 1482 184 1516
rect 218 1482 252 1516
rect 286 1482 345 1516
rect -11 1470 345 1482
<< psubdiffcont >>
rect 48 1482 82 1516
rect 116 1482 150 1516
rect 184 1482 218 1516
rect 252 1482 286 1516
<< poly >>
rect 0 1400 300 1430
rect 0 -48 300 0
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< polycont >>
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< locali >>
rect -9 1516 343 1526
rect -9 1482 42 1516
rect 82 1482 114 1516
rect 150 1482 184 1516
rect 220 1482 252 1516
rect 292 1482 343 1516
rect -9 1472 343 1482
rect 311 1363 345 1400
rect 311 1295 345 1329
rect 311 1227 345 1261
rect 311 1159 345 1193
rect 311 1091 345 1125
rect 311 1023 345 1057
rect 311 955 345 989
rect 311 887 345 921
rect 311 819 345 853
rect 311 751 345 785
rect 311 683 345 717
rect 311 615 345 649
rect 311 547 345 581
rect 311 479 345 513
rect 311 411 345 445
rect 311 343 345 377
rect 311 275 345 309
rect 311 207 345 241
rect 311 139 345 173
rect 311 71 345 105
rect 311 0 345 37
rect 0 -48 300 -42
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -88 300 -82
<< viali >>
rect 42 1482 48 1516
rect 48 1482 76 1516
rect 114 1482 116 1516
rect 116 1482 148 1516
rect 186 1482 218 1516
rect 218 1482 220 1516
rect 258 1482 286 1516
rect 286 1482 292 1516
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< metal1 >>
rect -9 1516 343 1526
rect -9 1482 42 1516
rect 76 1482 114 1516
rect 148 1482 186 1516
rect 220 1482 258 1516
rect 292 1482 343 1516
rect -9 1472 343 1482
rect 0 -48 300 -38
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< end >>
