magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 500
<< pwell >>
rect -37 -154 579 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -11 0 0 500
rect 500 471 553 500
rect 500 437 511 471
rect 545 437 553 471
rect 500 403 553 437
rect 500 369 511 403
rect 545 369 553 403
rect 500 335 553 369
rect 500 301 511 335
rect 545 301 553 335
rect 500 267 553 301
rect 500 233 511 267
rect 545 233 553 267
rect 500 199 553 233
rect 500 165 511 199
rect 545 165 553 199
rect 500 131 553 165
rect 500 97 511 131
rect 545 97 553 131
rect 500 63 553 97
rect 500 29 511 63
rect 545 29 553 63
rect 500 0 553 29
<< ndiffc >>
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< psubdiff >>
rect -11 -82 553 -70
rect -11 -116 16 -82
rect 50 -116 84 -82
rect 118 -116 152 -82
rect 186 -116 220 -82
rect 254 -116 288 -82
rect 322 -116 356 -82
rect 390 -116 424 -82
rect 458 -116 492 -82
rect 526 -116 553 -82
rect -11 -128 553 -116
<< psubdiffcont >>
rect 16 -116 50 -82
rect 84 -116 118 -82
rect 152 -116 186 -82
rect 220 -116 254 -82
rect 288 -116 322 -82
rect 356 -116 390 -82
rect 424 -116 458 -82
rect 492 -116 526 -82
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
rect -9 -82 551 -72
rect -9 -116 16 -82
rect 72 -116 84 -82
rect 144 -116 152 -82
rect 216 -116 220 -82
rect 322 -116 326 -82
rect 390 -116 398 -82
rect 458 -116 470 -82
rect 526 -116 551 -82
rect -9 -126 551 -116
<< viali >>
rect 38 -116 50 -82
rect 50 -116 72 -82
rect 110 -116 118 -82
rect 118 -116 144 -82
rect 182 -116 186 -82
rect 186 -116 216 -82
rect 254 -116 288 -82
rect 326 -116 356 -82
rect 356 -116 360 -82
rect 398 -116 424 -82
rect 424 -116 432 -82
rect 470 -116 492 -82
rect 492 -116 504 -82
<< metal1 >>
rect -9 -82 551 -72
rect -9 -116 38 -82
rect 72 -116 110 -82
rect 144 -116 182 -82
rect 216 -116 254 -82
rect 288 -116 326 -82
rect 360 -116 398 -82
rect 432 -116 470 -82
rect 504 -116 551 -82
rect -9 -126 551 -116
<< end >>
