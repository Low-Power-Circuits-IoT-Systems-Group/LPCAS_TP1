magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal3 >>
rect -2142 3787 -120 3820
rect -2142 3723 -204 3787
rect -140 3723 -120 3787
rect -2142 3707 -120 3723
rect -2142 3643 -204 3707
rect -140 3643 -120 3707
rect -2142 3627 -120 3643
rect -2142 3563 -204 3627
rect -140 3563 -120 3627
rect -2142 3547 -120 3563
rect -2142 3483 -204 3547
rect -140 3483 -120 3547
rect -2142 3467 -120 3483
rect -2142 3403 -204 3467
rect -140 3403 -120 3467
rect -2142 3387 -120 3403
rect -2142 3323 -204 3387
rect -140 3323 -120 3387
rect -2142 3307 -120 3323
rect -2142 3243 -204 3307
rect -140 3243 -120 3307
rect -2142 3227 -120 3243
rect -2142 3163 -204 3227
rect -140 3163 -120 3227
rect -2142 3147 -120 3163
rect -2142 3083 -204 3147
rect -140 3083 -120 3147
rect -2142 3067 -120 3083
rect -2142 3003 -204 3067
rect -140 3003 -120 3067
rect -2142 2987 -120 3003
rect -2142 2923 -204 2987
rect -140 2923 -120 2987
rect -2142 2907 -120 2923
rect -2142 2843 -204 2907
rect -140 2843 -120 2907
rect -2142 2827 -120 2843
rect -2142 2763 -204 2827
rect -140 2763 -120 2827
rect -2142 2747 -120 2763
rect -2142 2683 -204 2747
rect -140 2683 -120 2747
rect -2142 2667 -120 2683
rect -2142 2603 -204 2667
rect -140 2603 -120 2667
rect -2142 2587 -120 2603
rect -2142 2523 -204 2587
rect -140 2523 -120 2587
rect -2142 2507 -120 2523
rect -2142 2443 -204 2507
rect -140 2443 -120 2507
rect -2142 2427 -120 2443
rect -2142 2363 -204 2427
rect -140 2363 -120 2427
rect -2142 2347 -120 2363
rect -2142 2283 -204 2347
rect -140 2283 -120 2347
rect -2142 2267 -120 2283
rect -2142 2203 -204 2267
rect -140 2203 -120 2267
rect -2142 2187 -120 2203
rect -2142 2123 -204 2187
rect -140 2123 -120 2187
rect -2142 2090 -120 2123
rect 120 3787 2142 3820
rect 120 3723 2058 3787
rect 2122 3723 2142 3787
rect 120 3707 2142 3723
rect 120 3643 2058 3707
rect 2122 3643 2142 3707
rect 120 3627 2142 3643
rect 120 3563 2058 3627
rect 2122 3563 2142 3627
rect 120 3547 2142 3563
rect 120 3483 2058 3547
rect 2122 3483 2142 3547
rect 120 3467 2142 3483
rect 120 3403 2058 3467
rect 2122 3403 2142 3467
rect 120 3387 2142 3403
rect 120 3323 2058 3387
rect 2122 3323 2142 3387
rect 120 3307 2142 3323
rect 120 3243 2058 3307
rect 2122 3243 2142 3307
rect 120 3227 2142 3243
rect 120 3163 2058 3227
rect 2122 3163 2142 3227
rect 120 3147 2142 3163
rect 120 3083 2058 3147
rect 2122 3083 2142 3147
rect 120 3067 2142 3083
rect 120 3003 2058 3067
rect 2122 3003 2142 3067
rect 120 2987 2142 3003
rect 120 2923 2058 2987
rect 2122 2923 2142 2987
rect 120 2907 2142 2923
rect 120 2843 2058 2907
rect 2122 2843 2142 2907
rect 120 2827 2142 2843
rect 120 2763 2058 2827
rect 2122 2763 2142 2827
rect 120 2747 2142 2763
rect 120 2683 2058 2747
rect 2122 2683 2142 2747
rect 120 2667 2142 2683
rect 120 2603 2058 2667
rect 2122 2603 2142 2667
rect 120 2587 2142 2603
rect 120 2523 2058 2587
rect 2122 2523 2142 2587
rect 120 2507 2142 2523
rect 120 2443 2058 2507
rect 2122 2443 2142 2507
rect 120 2427 2142 2443
rect 120 2363 2058 2427
rect 2122 2363 2142 2427
rect 120 2347 2142 2363
rect 120 2283 2058 2347
rect 2122 2283 2142 2347
rect 120 2267 2142 2283
rect 120 2203 2058 2267
rect 2122 2203 2142 2267
rect 120 2187 2142 2203
rect 120 2123 2058 2187
rect 2122 2123 2142 2187
rect 120 2090 2142 2123
rect -2142 1817 -120 1850
rect -2142 1753 -204 1817
rect -140 1753 -120 1817
rect -2142 1737 -120 1753
rect -2142 1673 -204 1737
rect -140 1673 -120 1737
rect -2142 1657 -120 1673
rect -2142 1593 -204 1657
rect -140 1593 -120 1657
rect -2142 1577 -120 1593
rect -2142 1513 -204 1577
rect -140 1513 -120 1577
rect -2142 1497 -120 1513
rect -2142 1433 -204 1497
rect -140 1433 -120 1497
rect -2142 1417 -120 1433
rect -2142 1353 -204 1417
rect -140 1353 -120 1417
rect -2142 1337 -120 1353
rect -2142 1273 -204 1337
rect -140 1273 -120 1337
rect -2142 1257 -120 1273
rect -2142 1193 -204 1257
rect -140 1193 -120 1257
rect -2142 1177 -120 1193
rect -2142 1113 -204 1177
rect -140 1113 -120 1177
rect -2142 1097 -120 1113
rect -2142 1033 -204 1097
rect -140 1033 -120 1097
rect -2142 1017 -120 1033
rect -2142 953 -204 1017
rect -140 953 -120 1017
rect -2142 937 -120 953
rect -2142 873 -204 937
rect -140 873 -120 937
rect -2142 857 -120 873
rect -2142 793 -204 857
rect -140 793 -120 857
rect -2142 777 -120 793
rect -2142 713 -204 777
rect -140 713 -120 777
rect -2142 697 -120 713
rect -2142 633 -204 697
rect -140 633 -120 697
rect -2142 617 -120 633
rect -2142 553 -204 617
rect -140 553 -120 617
rect -2142 537 -120 553
rect -2142 473 -204 537
rect -140 473 -120 537
rect -2142 457 -120 473
rect -2142 393 -204 457
rect -140 393 -120 457
rect -2142 377 -120 393
rect -2142 313 -204 377
rect -140 313 -120 377
rect -2142 297 -120 313
rect -2142 233 -204 297
rect -140 233 -120 297
rect -2142 217 -120 233
rect -2142 153 -204 217
rect -140 153 -120 217
rect -2142 120 -120 153
rect 120 1817 2142 1850
rect 120 1753 2058 1817
rect 2122 1753 2142 1817
rect 120 1737 2142 1753
rect 120 1673 2058 1737
rect 2122 1673 2142 1737
rect 120 1657 2142 1673
rect 120 1593 2058 1657
rect 2122 1593 2142 1657
rect 120 1577 2142 1593
rect 120 1513 2058 1577
rect 2122 1513 2142 1577
rect 120 1497 2142 1513
rect 120 1433 2058 1497
rect 2122 1433 2142 1497
rect 120 1417 2142 1433
rect 120 1353 2058 1417
rect 2122 1353 2142 1417
rect 120 1337 2142 1353
rect 120 1273 2058 1337
rect 2122 1273 2142 1337
rect 120 1257 2142 1273
rect 120 1193 2058 1257
rect 2122 1193 2142 1257
rect 120 1177 2142 1193
rect 120 1113 2058 1177
rect 2122 1113 2142 1177
rect 120 1097 2142 1113
rect 120 1033 2058 1097
rect 2122 1033 2142 1097
rect 120 1017 2142 1033
rect 120 953 2058 1017
rect 2122 953 2142 1017
rect 120 937 2142 953
rect 120 873 2058 937
rect 2122 873 2142 937
rect 120 857 2142 873
rect 120 793 2058 857
rect 2122 793 2142 857
rect 120 777 2142 793
rect 120 713 2058 777
rect 2122 713 2142 777
rect 120 697 2142 713
rect 120 633 2058 697
rect 2122 633 2142 697
rect 120 617 2142 633
rect 120 553 2058 617
rect 2122 553 2142 617
rect 120 537 2142 553
rect 120 473 2058 537
rect 2122 473 2142 537
rect 120 457 2142 473
rect 120 393 2058 457
rect 2122 393 2142 457
rect 120 377 2142 393
rect 120 313 2058 377
rect 2122 313 2142 377
rect 120 297 2142 313
rect 120 233 2058 297
rect 2122 233 2142 297
rect 120 217 2142 233
rect 120 153 2058 217
rect 2122 153 2142 217
rect 120 120 2142 153
rect -2142 -153 -120 -120
rect -2142 -217 -204 -153
rect -140 -217 -120 -153
rect -2142 -233 -120 -217
rect -2142 -297 -204 -233
rect -140 -297 -120 -233
rect -2142 -313 -120 -297
rect -2142 -377 -204 -313
rect -140 -377 -120 -313
rect -2142 -393 -120 -377
rect -2142 -457 -204 -393
rect -140 -457 -120 -393
rect -2142 -473 -120 -457
rect -2142 -537 -204 -473
rect -140 -537 -120 -473
rect -2142 -553 -120 -537
rect -2142 -617 -204 -553
rect -140 -617 -120 -553
rect -2142 -633 -120 -617
rect -2142 -697 -204 -633
rect -140 -697 -120 -633
rect -2142 -713 -120 -697
rect -2142 -777 -204 -713
rect -140 -777 -120 -713
rect -2142 -793 -120 -777
rect -2142 -857 -204 -793
rect -140 -857 -120 -793
rect -2142 -873 -120 -857
rect -2142 -937 -204 -873
rect -140 -937 -120 -873
rect -2142 -953 -120 -937
rect -2142 -1017 -204 -953
rect -140 -1017 -120 -953
rect -2142 -1033 -120 -1017
rect -2142 -1097 -204 -1033
rect -140 -1097 -120 -1033
rect -2142 -1113 -120 -1097
rect -2142 -1177 -204 -1113
rect -140 -1177 -120 -1113
rect -2142 -1193 -120 -1177
rect -2142 -1257 -204 -1193
rect -140 -1257 -120 -1193
rect -2142 -1273 -120 -1257
rect -2142 -1337 -204 -1273
rect -140 -1337 -120 -1273
rect -2142 -1353 -120 -1337
rect -2142 -1417 -204 -1353
rect -140 -1417 -120 -1353
rect -2142 -1433 -120 -1417
rect -2142 -1497 -204 -1433
rect -140 -1497 -120 -1433
rect -2142 -1513 -120 -1497
rect -2142 -1577 -204 -1513
rect -140 -1577 -120 -1513
rect -2142 -1593 -120 -1577
rect -2142 -1657 -204 -1593
rect -140 -1657 -120 -1593
rect -2142 -1673 -120 -1657
rect -2142 -1737 -204 -1673
rect -140 -1737 -120 -1673
rect -2142 -1753 -120 -1737
rect -2142 -1817 -204 -1753
rect -140 -1817 -120 -1753
rect -2142 -1850 -120 -1817
rect 120 -153 2142 -120
rect 120 -217 2058 -153
rect 2122 -217 2142 -153
rect 120 -233 2142 -217
rect 120 -297 2058 -233
rect 2122 -297 2142 -233
rect 120 -313 2142 -297
rect 120 -377 2058 -313
rect 2122 -377 2142 -313
rect 120 -393 2142 -377
rect 120 -457 2058 -393
rect 2122 -457 2142 -393
rect 120 -473 2142 -457
rect 120 -537 2058 -473
rect 2122 -537 2142 -473
rect 120 -553 2142 -537
rect 120 -617 2058 -553
rect 2122 -617 2142 -553
rect 120 -633 2142 -617
rect 120 -697 2058 -633
rect 2122 -697 2142 -633
rect 120 -713 2142 -697
rect 120 -777 2058 -713
rect 2122 -777 2142 -713
rect 120 -793 2142 -777
rect 120 -857 2058 -793
rect 2122 -857 2142 -793
rect 120 -873 2142 -857
rect 120 -937 2058 -873
rect 2122 -937 2142 -873
rect 120 -953 2142 -937
rect 120 -1017 2058 -953
rect 2122 -1017 2142 -953
rect 120 -1033 2142 -1017
rect 120 -1097 2058 -1033
rect 2122 -1097 2142 -1033
rect 120 -1113 2142 -1097
rect 120 -1177 2058 -1113
rect 2122 -1177 2142 -1113
rect 120 -1193 2142 -1177
rect 120 -1257 2058 -1193
rect 2122 -1257 2142 -1193
rect 120 -1273 2142 -1257
rect 120 -1337 2058 -1273
rect 2122 -1337 2142 -1273
rect 120 -1353 2142 -1337
rect 120 -1417 2058 -1353
rect 2122 -1417 2142 -1353
rect 120 -1433 2142 -1417
rect 120 -1497 2058 -1433
rect 2122 -1497 2142 -1433
rect 120 -1513 2142 -1497
rect 120 -1577 2058 -1513
rect 2122 -1577 2142 -1513
rect 120 -1593 2142 -1577
rect 120 -1657 2058 -1593
rect 2122 -1657 2142 -1593
rect 120 -1673 2142 -1657
rect 120 -1737 2058 -1673
rect 2122 -1737 2142 -1673
rect 120 -1753 2142 -1737
rect 120 -1817 2058 -1753
rect 2122 -1817 2142 -1753
rect 120 -1850 2142 -1817
rect -2142 -2123 -120 -2090
rect -2142 -2187 -204 -2123
rect -140 -2187 -120 -2123
rect -2142 -2203 -120 -2187
rect -2142 -2267 -204 -2203
rect -140 -2267 -120 -2203
rect -2142 -2283 -120 -2267
rect -2142 -2347 -204 -2283
rect -140 -2347 -120 -2283
rect -2142 -2363 -120 -2347
rect -2142 -2427 -204 -2363
rect -140 -2427 -120 -2363
rect -2142 -2443 -120 -2427
rect -2142 -2507 -204 -2443
rect -140 -2507 -120 -2443
rect -2142 -2523 -120 -2507
rect -2142 -2587 -204 -2523
rect -140 -2587 -120 -2523
rect -2142 -2603 -120 -2587
rect -2142 -2667 -204 -2603
rect -140 -2667 -120 -2603
rect -2142 -2683 -120 -2667
rect -2142 -2747 -204 -2683
rect -140 -2747 -120 -2683
rect -2142 -2763 -120 -2747
rect -2142 -2827 -204 -2763
rect -140 -2827 -120 -2763
rect -2142 -2843 -120 -2827
rect -2142 -2907 -204 -2843
rect -140 -2907 -120 -2843
rect -2142 -2923 -120 -2907
rect -2142 -2987 -204 -2923
rect -140 -2987 -120 -2923
rect -2142 -3003 -120 -2987
rect -2142 -3067 -204 -3003
rect -140 -3067 -120 -3003
rect -2142 -3083 -120 -3067
rect -2142 -3147 -204 -3083
rect -140 -3147 -120 -3083
rect -2142 -3163 -120 -3147
rect -2142 -3227 -204 -3163
rect -140 -3227 -120 -3163
rect -2142 -3243 -120 -3227
rect -2142 -3307 -204 -3243
rect -140 -3307 -120 -3243
rect -2142 -3323 -120 -3307
rect -2142 -3387 -204 -3323
rect -140 -3387 -120 -3323
rect -2142 -3403 -120 -3387
rect -2142 -3467 -204 -3403
rect -140 -3467 -120 -3403
rect -2142 -3483 -120 -3467
rect -2142 -3547 -204 -3483
rect -140 -3547 -120 -3483
rect -2142 -3563 -120 -3547
rect -2142 -3627 -204 -3563
rect -140 -3627 -120 -3563
rect -2142 -3643 -120 -3627
rect -2142 -3707 -204 -3643
rect -140 -3707 -120 -3643
rect -2142 -3723 -120 -3707
rect -2142 -3787 -204 -3723
rect -140 -3787 -120 -3723
rect -2142 -3820 -120 -3787
rect 120 -2123 2142 -2090
rect 120 -2187 2058 -2123
rect 2122 -2187 2142 -2123
rect 120 -2203 2142 -2187
rect 120 -2267 2058 -2203
rect 2122 -2267 2142 -2203
rect 120 -2283 2142 -2267
rect 120 -2347 2058 -2283
rect 2122 -2347 2142 -2283
rect 120 -2363 2142 -2347
rect 120 -2427 2058 -2363
rect 2122 -2427 2142 -2363
rect 120 -2443 2142 -2427
rect 120 -2507 2058 -2443
rect 2122 -2507 2142 -2443
rect 120 -2523 2142 -2507
rect 120 -2587 2058 -2523
rect 2122 -2587 2142 -2523
rect 120 -2603 2142 -2587
rect 120 -2667 2058 -2603
rect 2122 -2667 2142 -2603
rect 120 -2683 2142 -2667
rect 120 -2747 2058 -2683
rect 2122 -2747 2142 -2683
rect 120 -2763 2142 -2747
rect 120 -2827 2058 -2763
rect 2122 -2827 2142 -2763
rect 120 -2843 2142 -2827
rect 120 -2907 2058 -2843
rect 2122 -2907 2142 -2843
rect 120 -2923 2142 -2907
rect 120 -2987 2058 -2923
rect 2122 -2987 2142 -2923
rect 120 -3003 2142 -2987
rect 120 -3067 2058 -3003
rect 2122 -3067 2142 -3003
rect 120 -3083 2142 -3067
rect 120 -3147 2058 -3083
rect 2122 -3147 2142 -3083
rect 120 -3163 2142 -3147
rect 120 -3227 2058 -3163
rect 2122 -3227 2142 -3163
rect 120 -3243 2142 -3227
rect 120 -3307 2058 -3243
rect 2122 -3307 2142 -3243
rect 120 -3323 2142 -3307
rect 120 -3387 2058 -3323
rect 2122 -3387 2142 -3323
rect 120 -3403 2142 -3387
rect 120 -3467 2058 -3403
rect 2122 -3467 2142 -3403
rect 120 -3483 2142 -3467
rect 120 -3547 2058 -3483
rect 2122 -3547 2142 -3483
rect 120 -3563 2142 -3547
rect 120 -3627 2058 -3563
rect 2122 -3627 2142 -3563
rect 120 -3643 2142 -3627
rect 120 -3707 2058 -3643
rect 2122 -3707 2142 -3643
rect 120 -3723 2142 -3707
rect 120 -3787 2058 -3723
rect 2122 -3787 2142 -3723
rect 120 -3820 2142 -3787
<< via3 >>
rect -204 3723 -140 3787
rect -204 3643 -140 3707
rect -204 3563 -140 3627
rect -204 3483 -140 3547
rect -204 3403 -140 3467
rect -204 3323 -140 3387
rect -204 3243 -140 3307
rect -204 3163 -140 3227
rect -204 3083 -140 3147
rect -204 3003 -140 3067
rect -204 2923 -140 2987
rect -204 2843 -140 2907
rect -204 2763 -140 2827
rect -204 2683 -140 2747
rect -204 2603 -140 2667
rect -204 2523 -140 2587
rect -204 2443 -140 2507
rect -204 2363 -140 2427
rect -204 2283 -140 2347
rect -204 2203 -140 2267
rect -204 2123 -140 2187
rect 2058 3723 2122 3787
rect 2058 3643 2122 3707
rect 2058 3563 2122 3627
rect 2058 3483 2122 3547
rect 2058 3403 2122 3467
rect 2058 3323 2122 3387
rect 2058 3243 2122 3307
rect 2058 3163 2122 3227
rect 2058 3083 2122 3147
rect 2058 3003 2122 3067
rect 2058 2923 2122 2987
rect 2058 2843 2122 2907
rect 2058 2763 2122 2827
rect 2058 2683 2122 2747
rect 2058 2603 2122 2667
rect 2058 2523 2122 2587
rect 2058 2443 2122 2507
rect 2058 2363 2122 2427
rect 2058 2283 2122 2347
rect 2058 2203 2122 2267
rect 2058 2123 2122 2187
rect -204 1753 -140 1817
rect -204 1673 -140 1737
rect -204 1593 -140 1657
rect -204 1513 -140 1577
rect -204 1433 -140 1497
rect -204 1353 -140 1417
rect -204 1273 -140 1337
rect -204 1193 -140 1257
rect -204 1113 -140 1177
rect -204 1033 -140 1097
rect -204 953 -140 1017
rect -204 873 -140 937
rect -204 793 -140 857
rect -204 713 -140 777
rect -204 633 -140 697
rect -204 553 -140 617
rect -204 473 -140 537
rect -204 393 -140 457
rect -204 313 -140 377
rect -204 233 -140 297
rect -204 153 -140 217
rect 2058 1753 2122 1817
rect 2058 1673 2122 1737
rect 2058 1593 2122 1657
rect 2058 1513 2122 1577
rect 2058 1433 2122 1497
rect 2058 1353 2122 1417
rect 2058 1273 2122 1337
rect 2058 1193 2122 1257
rect 2058 1113 2122 1177
rect 2058 1033 2122 1097
rect 2058 953 2122 1017
rect 2058 873 2122 937
rect 2058 793 2122 857
rect 2058 713 2122 777
rect 2058 633 2122 697
rect 2058 553 2122 617
rect 2058 473 2122 537
rect 2058 393 2122 457
rect 2058 313 2122 377
rect 2058 233 2122 297
rect 2058 153 2122 217
rect -204 -217 -140 -153
rect -204 -297 -140 -233
rect -204 -377 -140 -313
rect -204 -457 -140 -393
rect -204 -537 -140 -473
rect -204 -617 -140 -553
rect -204 -697 -140 -633
rect -204 -777 -140 -713
rect -204 -857 -140 -793
rect -204 -937 -140 -873
rect -204 -1017 -140 -953
rect -204 -1097 -140 -1033
rect -204 -1177 -140 -1113
rect -204 -1257 -140 -1193
rect -204 -1337 -140 -1273
rect -204 -1417 -140 -1353
rect -204 -1497 -140 -1433
rect -204 -1577 -140 -1513
rect -204 -1657 -140 -1593
rect -204 -1737 -140 -1673
rect -204 -1817 -140 -1753
rect 2058 -217 2122 -153
rect 2058 -297 2122 -233
rect 2058 -377 2122 -313
rect 2058 -457 2122 -393
rect 2058 -537 2122 -473
rect 2058 -617 2122 -553
rect 2058 -697 2122 -633
rect 2058 -777 2122 -713
rect 2058 -857 2122 -793
rect 2058 -937 2122 -873
rect 2058 -1017 2122 -953
rect 2058 -1097 2122 -1033
rect 2058 -1177 2122 -1113
rect 2058 -1257 2122 -1193
rect 2058 -1337 2122 -1273
rect 2058 -1417 2122 -1353
rect 2058 -1497 2122 -1433
rect 2058 -1577 2122 -1513
rect 2058 -1657 2122 -1593
rect 2058 -1737 2122 -1673
rect 2058 -1817 2122 -1753
rect -204 -2187 -140 -2123
rect -204 -2267 -140 -2203
rect -204 -2347 -140 -2283
rect -204 -2427 -140 -2363
rect -204 -2507 -140 -2443
rect -204 -2587 -140 -2523
rect -204 -2667 -140 -2603
rect -204 -2747 -140 -2683
rect -204 -2827 -140 -2763
rect -204 -2907 -140 -2843
rect -204 -2987 -140 -2923
rect -204 -3067 -140 -3003
rect -204 -3147 -140 -3083
rect -204 -3227 -140 -3163
rect -204 -3307 -140 -3243
rect -204 -3387 -140 -3323
rect -204 -3467 -140 -3403
rect -204 -3547 -140 -3483
rect -204 -3627 -140 -3563
rect -204 -3707 -140 -3643
rect -204 -3787 -140 -3723
rect 2058 -2187 2122 -2123
rect 2058 -2267 2122 -2203
rect 2058 -2347 2122 -2283
rect 2058 -2427 2122 -2363
rect 2058 -2507 2122 -2443
rect 2058 -2587 2122 -2523
rect 2058 -2667 2122 -2603
rect 2058 -2747 2122 -2683
rect 2058 -2827 2122 -2763
rect 2058 -2907 2122 -2843
rect 2058 -2987 2122 -2923
rect 2058 -3067 2122 -3003
rect 2058 -3147 2122 -3083
rect 2058 -3227 2122 -3163
rect 2058 -3307 2122 -3243
rect 2058 -3387 2122 -3323
rect 2058 -3467 2122 -3403
rect 2058 -3547 2122 -3483
rect 2058 -3627 2122 -3563
rect 2058 -3707 2122 -3643
rect 2058 -3787 2122 -3723
<< mimcap >>
rect -2102 3707 -452 3780
rect -2102 2203 -2029 3707
rect -525 2203 -452 3707
rect -2102 2130 -452 2203
rect 160 3707 1810 3780
rect 160 2203 233 3707
rect 1737 2203 1810 3707
rect 160 2130 1810 2203
rect -2102 1737 -452 1810
rect -2102 233 -2029 1737
rect -525 233 -452 1737
rect -2102 160 -452 233
rect 160 1737 1810 1810
rect 160 233 233 1737
rect 1737 233 1810 1737
rect 160 160 1810 233
rect -2102 -233 -452 -160
rect -2102 -1737 -2029 -233
rect -525 -1737 -452 -233
rect -2102 -1810 -452 -1737
rect 160 -233 1810 -160
rect 160 -1737 233 -233
rect 1737 -1737 1810 -233
rect 160 -1810 1810 -1737
rect -2102 -2203 -452 -2130
rect -2102 -3707 -2029 -2203
rect -525 -3707 -452 -2203
rect -2102 -3780 -452 -3707
rect 160 -2203 1810 -2130
rect 160 -3707 233 -2203
rect 1737 -3707 1810 -2203
rect 160 -3780 1810 -3707
<< mimcapcontact >>
rect -2029 2203 -525 3707
rect 233 2203 1737 3707
rect -2029 233 -525 1737
rect 233 233 1737 1737
rect -2029 -1737 -525 -233
rect 233 -1737 1737 -233
rect -2029 -3707 -525 -2203
rect 233 -3707 1737 -2203
<< metal4 >>
rect -1329 3741 -1225 3940
rect -224 3787 -120 3940
rect -2063 3707 -491 3741
rect -2063 2203 -2029 3707
rect -525 2203 -491 3707
rect -2063 2169 -491 2203
rect -224 3723 -204 3787
rect -140 3723 -120 3787
rect 933 3741 1037 3940
rect 2038 3787 2142 3940
rect -224 3707 -120 3723
rect -224 3643 -204 3707
rect -140 3643 -120 3707
rect -224 3627 -120 3643
rect -224 3563 -204 3627
rect -140 3563 -120 3627
rect -224 3547 -120 3563
rect -224 3483 -204 3547
rect -140 3483 -120 3547
rect -224 3467 -120 3483
rect -224 3403 -204 3467
rect -140 3403 -120 3467
rect -224 3387 -120 3403
rect -224 3323 -204 3387
rect -140 3323 -120 3387
rect -224 3307 -120 3323
rect -224 3243 -204 3307
rect -140 3243 -120 3307
rect -224 3227 -120 3243
rect -224 3163 -204 3227
rect -140 3163 -120 3227
rect -224 3147 -120 3163
rect -224 3083 -204 3147
rect -140 3083 -120 3147
rect -224 3067 -120 3083
rect -224 3003 -204 3067
rect -140 3003 -120 3067
rect -224 2987 -120 3003
rect -224 2923 -204 2987
rect -140 2923 -120 2987
rect -224 2907 -120 2923
rect -224 2843 -204 2907
rect -140 2843 -120 2907
rect -224 2827 -120 2843
rect -224 2763 -204 2827
rect -140 2763 -120 2827
rect -224 2747 -120 2763
rect -224 2683 -204 2747
rect -140 2683 -120 2747
rect -224 2667 -120 2683
rect -224 2603 -204 2667
rect -140 2603 -120 2667
rect -224 2587 -120 2603
rect -224 2523 -204 2587
rect -140 2523 -120 2587
rect -224 2507 -120 2523
rect -224 2443 -204 2507
rect -140 2443 -120 2507
rect -224 2427 -120 2443
rect -224 2363 -204 2427
rect -140 2363 -120 2427
rect -224 2347 -120 2363
rect -224 2283 -204 2347
rect -140 2283 -120 2347
rect -224 2267 -120 2283
rect -224 2203 -204 2267
rect -140 2203 -120 2267
rect -224 2187 -120 2203
rect -1329 1771 -1225 2169
rect -224 2123 -204 2187
rect -140 2123 -120 2187
rect 199 3707 1771 3741
rect 199 2203 233 3707
rect 1737 2203 1771 3707
rect 199 2169 1771 2203
rect 2038 3723 2058 3787
rect 2122 3723 2142 3787
rect 2038 3707 2142 3723
rect 2038 3643 2058 3707
rect 2122 3643 2142 3707
rect 2038 3627 2142 3643
rect 2038 3563 2058 3627
rect 2122 3563 2142 3627
rect 2038 3547 2142 3563
rect 2038 3483 2058 3547
rect 2122 3483 2142 3547
rect 2038 3467 2142 3483
rect 2038 3403 2058 3467
rect 2122 3403 2142 3467
rect 2038 3387 2142 3403
rect 2038 3323 2058 3387
rect 2122 3323 2142 3387
rect 2038 3307 2142 3323
rect 2038 3243 2058 3307
rect 2122 3243 2142 3307
rect 2038 3227 2142 3243
rect 2038 3163 2058 3227
rect 2122 3163 2142 3227
rect 2038 3147 2142 3163
rect 2038 3083 2058 3147
rect 2122 3083 2142 3147
rect 2038 3067 2142 3083
rect 2038 3003 2058 3067
rect 2122 3003 2142 3067
rect 2038 2987 2142 3003
rect 2038 2923 2058 2987
rect 2122 2923 2142 2987
rect 2038 2907 2142 2923
rect 2038 2843 2058 2907
rect 2122 2843 2142 2907
rect 2038 2827 2142 2843
rect 2038 2763 2058 2827
rect 2122 2763 2142 2827
rect 2038 2747 2142 2763
rect 2038 2683 2058 2747
rect 2122 2683 2142 2747
rect 2038 2667 2142 2683
rect 2038 2603 2058 2667
rect 2122 2603 2142 2667
rect 2038 2587 2142 2603
rect 2038 2523 2058 2587
rect 2122 2523 2142 2587
rect 2038 2507 2142 2523
rect 2038 2443 2058 2507
rect 2122 2443 2142 2507
rect 2038 2427 2142 2443
rect 2038 2363 2058 2427
rect 2122 2363 2142 2427
rect 2038 2347 2142 2363
rect 2038 2283 2058 2347
rect 2122 2283 2142 2347
rect 2038 2267 2142 2283
rect 2038 2203 2058 2267
rect 2122 2203 2142 2267
rect 2038 2187 2142 2203
rect -224 1817 -120 2123
rect -2063 1737 -491 1771
rect -2063 233 -2029 1737
rect -525 233 -491 1737
rect -2063 199 -491 233
rect -224 1753 -204 1817
rect -140 1753 -120 1817
rect 933 1771 1037 2169
rect 2038 2123 2058 2187
rect 2122 2123 2142 2187
rect 2038 1817 2142 2123
rect -224 1737 -120 1753
rect -224 1673 -204 1737
rect -140 1673 -120 1737
rect -224 1657 -120 1673
rect -224 1593 -204 1657
rect -140 1593 -120 1657
rect -224 1577 -120 1593
rect -224 1513 -204 1577
rect -140 1513 -120 1577
rect -224 1497 -120 1513
rect -224 1433 -204 1497
rect -140 1433 -120 1497
rect -224 1417 -120 1433
rect -224 1353 -204 1417
rect -140 1353 -120 1417
rect -224 1337 -120 1353
rect -224 1273 -204 1337
rect -140 1273 -120 1337
rect -224 1257 -120 1273
rect -224 1193 -204 1257
rect -140 1193 -120 1257
rect -224 1177 -120 1193
rect -224 1113 -204 1177
rect -140 1113 -120 1177
rect -224 1097 -120 1113
rect -224 1033 -204 1097
rect -140 1033 -120 1097
rect -224 1017 -120 1033
rect -224 953 -204 1017
rect -140 953 -120 1017
rect -224 937 -120 953
rect -224 873 -204 937
rect -140 873 -120 937
rect -224 857 -120 873
rect -224 793 -204 857
rect -140 793 -120 857
rect -224 777 -120 793
rect -224 713 -204 777
rect -140 713 -120 777
rect -224 697 -120 713
rect -224 633 -204 697
rect -140 633 -120 697
rect -224 617 -120 633
rect -224 553 -204 617
rect -140 553 -120 617
rect -224 537 -120 553
rect -224 473 -204 537
rect -140 473 -120 537
rect -224 457 -120 473
rect -224 393 -204 457
rect -140 393 -120 457
rect -224 377 -120 393
rect -224 313 -204 377
rect -140 313 -120 377
rect -224 297 -120 313
rect -224 233 -204 297
rect -140 233 -120 297
rect -224 217 -120 233
rect -1329 -199 -1225 199
rect -224 153 -204 217
rect -140 153 -120 217
rect 199 1737 1771 1771
rect 199 233 233 1737
rect 1737 233 1771 1737
rect 199 199 1771 233
rect 2038 1753 2058 1817
rect 2122 1753 2142 1817
rect 2038 1737 2142 1753
rect 2038 1673 2058 1737
rect 2122 1673 2142 1737
rect 2038 1657 2142 1673
rect 2038 1593 2058 1657
rect 2122 1593 2142 1657
rect 2038 1577 2142 1593
rect 2038 1513 2058 1577
rect 2122 1513 2142 1577
rect 2038 1497 2142 1513
rect 2038 1433 2058 1497
rect 2122 1433 2142 1497
rect 2038 1417 2142 1433
rect 2038 1353 2058 1417
rect 2122 1353 2142 1417
rect 2038 1337 2142 1353
rect 2038 1273 2058 1337
rect 2122 1273 2142 1337
rect 2038 1257 2142 1273
rect 2038 1193 2058 1257
rect 2122 1193 2142 1257
rect 2038 1177 2142 1193
rect 2038 1113 2058 1177
rect 2122 1113 2142 1177
rect 2038 1097 2142 1113
rect 2038 1033 2058 1097
rect 2122 1033 2142 1097
rect 2038 1017 2142 1033
rect 2038 953 2058 1017
rect 2122 953 2142 1017
rect 2038 937 2142 953
rect 2038 873 2058 937
rect 2122 873 2142 937
rect 2038 857 2142 873
rect 2038 793 2058 857
rect 2122 793 2142 857
rect 2038 777 2142 793
rect 2038 713 2058 777
rect 2122 713 2142 777
rect 2038 697 2142 713
rect 2038 633 2058 697
rect 2122 633 2142 697
rect 2038 617 2142 633
rect 2038 553 2058 617
rect 2122 553 2142 617
rect 2038 537 2142 553
rect 2038 473 2058 537
rect 2122 473 2142 537
rect 2038 457 2142 473
rect 2038 393 2058 457
rect 2122 393 2142 457
rect 2038 377 2142 393
rect 2038 313 2058 377
rect 2122 313 2142 377
rect 2038 297 2142 313
rect 2038 233 2058 297
rect 2122 233 2142 297
rect 2038 217 2142 233
rect -224 -153 -120 153
rect -2063 -233 -491 -199
rect -2063 -1737 -2029 -233
rect -525 -1737 -491 -233
rect -2063 -1771 -491 -1737
rect -224 -217 -204 -153
rect -140 -217 -120 -153
rect 933 -199 1037 199
rect 2038 153 2058 217
rect 2122 153 2142 217
rect 2038 -153 2142 153
rect -224 -233 -120 -217
rect -224 -297 -204 -233
rect -140 -297 -120 -233
rect -224 -313 -120 -297
rect -224 -377 -204 -313
rect -140 -377 -120 -313
rect -224 -393 -120 -377
rect -224 -457 -204 -393
rect -140 -457 -120 -393
rect -224 -473 -120 -457
rect -224 -537 -204 -473
rect -140 -537 -120 -473
rect -224 -553 -120 -537
rect -224 -617 -204 -553
rect -140 -617 -120 -553
rect -224 -633 -120 -617
rect -224 -697 -204 -633
rect -140 -697 -120 -633
rect -224 -713 -120 -697
rect -224 -777 -204 -713
rect -140 -777 -120 -713
rect -224 -793 -120 -777
rect -224 -857 -204 -793
rect -140 -857 -120 -793
rect -224 -873 -120 -857
rect -224 -937 -204 -873
rect -140 -937 -120 -873
rect -224 -953 -120 -937
rect -224 -1017 -204 -953
rect -140 -1017 -120 -953
rect -224 -1033 -120 -1017
rect -224 -1097 -204 -1033
rect -140 -1097 -120 -1033
rect -224 -1113 -120 -1097
rect -224 -1177 -204 -1113
rect -140 -1177 -120 -1113
rect -224 -1193 -120 -1177
rect -224 -1257 -204 -1193
rect -140 -1257 -120 -1193
rect -224 -1273 -120 -1257
rect -224 -1337 -204 -1273
rect -140 -1337 -120 -1273
rect -224 -1353 -120 -1337
rect -224 -1417 -204 -1353
rect -140 -1417 -120 -1353
rect -224 -1433 -120 -1417
rect -224 -1497 -204 -1433
rect -140 -1497 -120 -1433
rect -224 -1513 -120 -1497
rect -224 -1577 -204 -1513
rect -140 -1577 -120 -1513
rect -224 -1593 -120 -1577
rect -224 -1657 -204 -1593
rect -140 -1657 -120 -1593
rect -224 -1673 -120 -1657
rect -224 -1737 -204 -1673
rect -140 -1737 -120 -1673
rect -224 -1753 -120 -1737
rect -1329 -2169 -1225 -1771
rect -224 -1817 -204 -1753
rect -140 -1817 -120 -1753
rect 199 -233 1771 -199
rect 199 -1737 233 -233
rect 1737 -1737 1771 -233
rect 199 -1771 1771 -1737
rect 2038 -217 2058 -153
rect 2122 -217 2142 -153
rect 2038 -233 2142 -217
rect 2038 -297 2058 -233
rect 2122 -297 2142 -233
rect 2038 -313 2142 -297
rect 2038 -377 2058 -313
rect 2122 -377 2142 -313
rect 2038 -393 2142 -377
rect 2038 -457 2058 -393
rect 2122 -457 2142 -393
rect 2038 -473 2142 -457
rect 2038 -537 2058 -473
rect 2122 -537 2142 -473
rect 2038 -553 2142 -537
rect 2038 -617 2058 -553
rect 2122 -617 2142 -553
rect 2038 -633 2142 -617
rect 2038 -697 2058 -633
rect 2122 -697 2142 -633
rect 2038 -713 2142 -697
rect 2038 -777 2058 -713
rect 2122 -777 2142 -713
rect 2038 -793 2142 -777
rect 2038 -857 2058 -793
rect 2122 -857 2142 -793
rect 2038 -873 2142 -857
rect 2038 -937 2058 -873
rect 2122 -937 2142 -873
rect 2038 -953 2142 -937
rect 2038 -1017 2058 -953
rect 2122 -1017 2142 -953
rect 2038 -1033 2142 -1017
rect 2038 -1097 2058 -1033
rect 2122 -1097 2142 -1033
rect 2038 -1113 2142 -1097
rect 2038 -1177 2058 -1113
rect 2122 -1177 2142 -1113
rect 2038 -1193 2142 -1177
rect 2038 -1257 2058 -1193
rect 2122 -1257 2142 -1193
rect 2038 -1273 2142 -1257
rect 2038 -1337 2058 -1273
rect 2122 -1337 2142 -1273
rect 2038 -1353 2142 -1337
rect 2038 -1417 2058 -1353
rect 2122 -1417 2142 -1353
rect 2038 -1433 2142 -1417
rect 2038 -1497 2058 -1433
rect 2122 -1497 2142 -1433
rect 2038 -1513 2142 -1497
rect 2038 -1577 2058 -1513
rect 2122 -1577 2142 -1513
rect 2038 -1593 2142 -1577
rect 2038 -1657 2058 -1593
rect 2122 -1657 2142 -1593
rect 2038 -1673 2142 -1657
rect 2038 -1737 2058 -1673
rect 2122 -1737 2142 -1673
rect 2038 -1753 2142 -1737
rect -224 -2123 -120 -1817
rect -2063 -2203 -491 -2169
rect -2063 -3707 -2029 -2203
rect -525 -3707 -491 -2203
rect -2063 -3741 -491 -3707
rect -224 -2187 -204 -2123
rect -140 -2187 -120 -2123
rect 933 -2169 1037 -1771
rect 2038 -1817 2058 -1753
rect 2122 -1817 2142 -1753
rect 2038 -2123 2142 -1817
rect -224 -2203 -120 -2187
rect -224 -2267 -204 -2203
rect -140 -2267 -120 -2203
rect -224 -2283 -120 -2267
rect -224 -2347 -204 -2283
rect -140 -2347 -120 -2283
rect -224 -2363 -120 -2347
rect -224 -2427 -204 -2363
rect -140 -2427 -120 -2363
rect -224 -2443 -120 -2427
rect -224 -2507 -204 -2443
rect -140 -2507 -120 -2443
rect -224 -2523 -120 -2507
rect -224 -2587 -204 -2523
rect -140 -2587 -120 -2523
rect -224 -2603 -120 -2587
rect -224 -2667 -204 -2603
rect -140 -2667 -120 -2603
rect -224 -2683 -120 -2667
rect -224 -2747 -204 -2683
rect -140 -2747 -120 -2683
rect -224 -2763 -120 -2747
rect -224 -2827 -204 -2763
rect -140 -2827 -120 -2763
rect -224 -2843 -120 -2827
rect -224 -2907 -204 -2843
rect -140 -2907 -120 -2843
rect -224 -2923 -120 -2907
rect -224 -2987 -204 -2923
rect -140 -2987 -120 -2923
rect -224 -3003 -120 -2987
rect -224 -3067 -204 -3003
rect -140 -3067 -120 -3003
rect -224 -3083 -120 -3067
rect -224 -3147 -204 -3083
rect -140 -3147 -120 -3083
rect -224 -3163 -120 -3147
rect -224 -3227 -204 -3163
rect -140 -3227 -120 -3163
rect -224 -3243 -120 -3227
rect -224 -3307 -204 -3243
rect -140 -3307 -120 -3243
rect -224 -3323 -120 -3307
rect -224 -3387 -204 -3323
rect -140 -3387 -120 -3323
rect -224 -3403 -120 -3387
rect -224 -3467 -204 -3403
rect -140 -3467 -120 -3403
rect -224 -3483 -120 -3467
rect -224 -3547 -204 -3483
rect -140 -3547 -120 -3483
rect -224 -3563 -120 -3547
rect -224 -3627 -204 -3563
rect -140 -3627 -120 -3563
rect -224 -3643 -120 -3627
rect -224 -3707 -204 -3643
rect -140 -3707 -120 -3643
rect -224 -3723 -120 -3707
rect -1329 -3940 -1225 -3741
rect -224 -3787 -204 -3723
rect -140 -3787 -120 -3723
rect 199 -2203 1771 -2169
rect 199 -3707 233 -2203
rect 1737 -3707 1771 -2203
rect 199 -3741 1771 -3707
rect 2038 -2187 2058 -2123
rect 2122 -2187 2142 -2123
rect 2038 -2203 2142 -2187
rect 2038 -2267 2058 -2203
rect 2122 -2267 2142 -2203
rect 2038 -2283 2142 -2267
rect 2038 -2347 2058 -2283
rect 2122 -2347 2142 -2283
rect 2038 -2363 2142 -2347
rect 2038 -2427 2058 -2363
rect 2122 -2427 2142 -2363
rect 2038 -2443 2142 -2427
rect 2038 -2507 2058 -2443
rect 2122 -2507 2142 -2443
rect 2038 -2523 2142 -2507
rect 2038 -2587 2058 -2523
rect 2122 -2587 2142 -2523
rect 2038 -2603 2142 -2587
rect 2038 -2667 2058 -2603
rect 2122 -2667 2142 -2603
rect 2038 -2683 2142 -2667
rect 2038 -2747 2058 -2683
rect 2122 -2747 2142 -2683
rect 2038 -2763 2142 -2747
rect 2038 -2827 2058 -2763
rect 2122 -2827 2142 -2763
rect 2038 -2843 2142 -2827
rect 2038 -2907 2058 -2843
rect 2122 -2907 2142 -2843
rect 2038 -2923 2142 -2907
rect 2038 -2987 2058 -2923
rect 2122 -2987 2142 -2923
rect 2038 -3003 2142 -2987
rect 2038 -3067 2058 -3003
rect 2122 -3067 2142 -3003
rect 2038 -3083 2142 -3067
rect 2038 -3147 2058 -3083
rect 2122 -3147 2142 -3083
rect 2038 -3163 2142 -3147
rect 2038 -3227 2058 -3163
rect 2122 -3227 2142 -3163
rect 2038 -3243 2142 -3227
rect 2038 -3307 2058 -3243
rect 2122 -3307 2142 -3243
rect 2038 -3323 2142 -3307
rect 2038 -3387 2058 -3323
rect 2122 -3387 2142 -3323
rect 2038 -3403 2142 -3387
rect 2038 -3467 2058 -3403
rect 2122 -3467 2142 -3403
rect 2038 -3483 2142 -3467
rect 2038 -3547 2058 -3483
rect 2122 -3547 2142 -3483
rect 2038 -3563 2142 -3547
rect 2038 -3627 2058 -3563
rect 2122 -3627 2142 -3563
rect 2038 -3643 2142 -3627
rect 2038 -3707 2058 -3643
rect 2122 -3707 2142 -3643
rect 2038 -3723 2142 -3707
rect -224 -3940 -120 -3787
rect 933 -3940 1037 -3741
rect 2038 -3787 2058 -3723
rect 2122 -3787 2142 -3723
rect 2038 -3940 2142 -3787
<< properties >>
string FIXED_BBOX 120 2090 1850 3820
<< end >>
