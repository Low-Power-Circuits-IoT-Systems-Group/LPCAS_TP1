magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 600
rect 245 555 250 600
rect 237 521 250 555
rect 245 487 250 521
rect 237 453 250 487
rect 245 419 250 453
rect 237 385 250 419
rect 245 351 250 385
rect 237 317 250 351
rect 245 283 250 317
rect 237 249 250 283
rect 245 215 250 249
rect 237 181 250 215
rect 245 147 250 181
rect 237 113 250 147
rect 245 79 250 113
rect 237 45 250 79
rect 245 0 250 45
<< nwell >>
rect -47 -36 281 636
<< pmos >>
rect 0 0 200 600
<< pdiff >>
rect -11 0 0 600
rect 200 555 245 600
rect 200 521 211 555
rect 200 487 245 521
rect 200 453 211 487
rect 200 419 245 453
rect 200 385 211 419
rect 200 351 245 385
rect 200 317 211 351
rect 200 283 245 317
rect 200 249 211 283
rect 200 215 245 249
rect 200 181 211 215
rect 200 147 245 181
rect 200 113 211 147
rect 200 79 245 113
rect 200 45 211 79
rect 200 0 245 45
<< pdiffc >>
rect 211 521 245 555
rect 211 453 245 487
rect 211 385 245 419
rect 211 317 245 351
rect 211 249 245 283
rect 211 181 245 215
rect 211 113 245 147
rect 211 45 245 79
<< poly >>
rect 0 682 200 692
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 600 200 648
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 648 50 682
rect 150 648 184 682
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect 0 682 200 688
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 642 200 648
rect 211 555 245 600
rect 211 487 245 521
rect 211 419 245 453
rect 211 351 245 385
rect 211 283 245 317
rect 211 215 245 249
rect 211 147 245 181
rect 211 79 245 113
rect 211 0 245 45
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect 16 648 50 682
rect 150 648 184 682
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect 0 682 200 692
rect 0 648 16 682
rect 50 648 150 682
rect 184 648 200 682
rect 0 638 200 648
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
