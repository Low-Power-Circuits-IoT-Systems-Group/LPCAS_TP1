magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 2000
rect 75 1969 80 2000
rect 67 1935 80 1969
rect 75 1901 80 1935
rect 67 1867 80 1901
rect 75 1833 80 1867
rect 67 1799 80 1833
rect 75 1765 80 1799
rect 67 1731 80 1765
rect 75 1697 80 1731
rect 67 1663 80 1697
rect 75 1629 80 1663
rect 67 1595 80 1629
rect 75 1561 80 1595
rect 67 1527 80 1561
rect 75 1493 80 1527
rect 67 1459 80 1493
rect 75 1425 80 1459
rect 67 1391 80 1425
rect 75 1357 80 1391
rect 67 1323 80 1357
rect 75 1289 80 1323
rect 67 1255 80 1289
rect 75 1221 80 1255
rect 67 1187 80 1221
rect 75 1153 80 1187
rect 67 1119 80 1153
rect 75 1085 80 1119
rect 67 1051 80 1085
rect 75 1017 80 1051
rect 67 983 80 1017
rect 75 949 80 983
rect 67 915 80 949
rect 75 881 80 915
rect 67 847 80 881
rect 75 813 80 847
rect 67 779 80 813
rect 75 745 80 779
rect 67 711 80 745
rect 75 677 80 711
rect 67 643 80 677
rect 75 609 80 643
rect 67 575 80 609
rect 75 541 80 575
rect 67 507 80 541
rect 75 473 80 507
rect 67 439 80 473
rect 75 405 80 439
rect 67 371 80 405
rect 75 337 80 371
rect 67 303 80 337
rect 75 269 80 303
rect 67 235 80 269
rect 75 201 80 235
rect 67 167 80 201
rect 75 133 80 167
rect 67 99 80 133
rect 75 65 80 99
rect 67 31 80 65
rect 75 0 80 31
<< pwell >>
rect -37 -154 101 2026
<< nmos >>
rect 0 0 30 2000
<< ndiff >>
rect -11 0 0 2000
rect 30 1969 75 2000
rect 30 1935 41 1969
rect 30 1901 75 1935
rect 30 1867 41 1901
rect 30 1833 75 1867
rect 30 1799 41 1833
rect 30 1765 75 1799
rect 30 1731 41 1765
rect 30 1697 75 1731
rect 30 1663 41 1697
rect 30 1629 75 1663
rect 30 1595 41 1629
rect 30 1561 75 1595
rect 30 1527 41 1561
rect 30 1493 75 1527
rect 30 1459 41 1493
rect 30 1425 75 1459
rect 30 1391 41 1425
rect 30 1357 75 1391
rect 30 1323 41 1357
rect 30 1289 75 1323
rect 30 1255 41 1289
rect 30 1221 75 1255
rect 30 1187 41 1221
rect 30 1153 75 1187
rect 30 1119 41 1153
rect 30 1085 75 1119
rect 30 1051 41 1085
rect 30 1017 75 1051
rect 30 983 41 1017
rect 30 949 75 983
rect 30 915 41 949
rect 30 881 75 915
rect 30 847 41 881
rect 30 813 75 847
rect 30 779 41 813
rect 30 745 75 779
rect 30 711 41 745
rect 30 677 75 711
rect 30 643 41 677
rect 30 609 75 643
rect 30 575 41 609
rect 30 541 75 575
rect 30 507 41 541
rect 30 473 75 507
rect 30 439 41 473
rect 30 405 75 439
rect 30 371 41 405
rect 30 337 75 371
rect 30 303 41 337
rect 30 269 75 303
rect 30 235 41 269
rect 30 201 75 235
rect 30 167 41 201
rect 30 133 75 167
rect 30 99 41 133
rect 30 65 75 99
rect 30 31 41 65
rect 30 0 75 31
<< ndiffc >>
rect 41 1935 75 1969
rect 41 1867 75 1901
rect 41 1799 75 1833
rect 41 1731 75 1765
rect 41 1663 75 1697
rect 41 1595 75 1629
rect 41 1527 75 1561
rect 41 1459 75 1493
rect 41 1391 75 1425
rect 41 1323 75 1357
rect 41 1255 75 1289
rect 41 1187 75 1221
rect 41 1119 75 1153
rect 41 1051 75 1085
rect 41 983 75 1017
rect 41 915 75 949
rect 41 847 75 881
rect 41 779 75 813
rect 41 711 75 745
rect 41 643 75 677
rect 41 575 75 609
rect 41 507 75 541
rect 41 439 75 473
rect 41 371 75 405
rect 41 303 75 337
rect 41 235 75 269
rect 41 167 75 201
rect 41 99 75 133
rect 41 31 75 65
<< psubdiff >>
rect -11 -82 75 -70
rect -11 -116 15 -82
rect 49 -116 75 -82
rect -11 -128 75 -116
<< psubdiffcont >>
rect 15 -116 49 -82
<< poly >>
rect 0 2000 30 2030
rect 0 -30 30 0
<< locali >>
rect 41 1969 75 2000
rect 41 1901 75 1935
rect 41 1833 75 1867
rect 41 1765 75 1799
rect 41 1697 75 1731
rect 41 1629 75 1663
rect 41 1561 75 1595
rect 41 1493 75 1527
rect 41 1425 75 1459
rect 41 1357 75 1391
rect 41 1289 75 1323
rect 41 1221 75 1255
rect 41 1153 75 1187
rect 41 1085 75 1119
rect 41 1017 75 1051
rect 41 949 75 983
rect 41 881 75 915
rect 41 813 75 847
rect 41 745 75 779
rect 41 677 75 711
rect 41 609 75 643
rect 41 541 75 575
rect 41 473 75 507
rect 41 405 75 439
rect 41 337 75 371
rect 41 269 75 303
rect 41 201 75 235
rect 41 133 75 167
rect 41 65 75 99
rect 41 0 75 31
rect -9 -82 73 -72
rect -9 -116 15 -82
rect 49 -116 73 -82
rect -9 -126 73 -116
<< viali >>
rect 15 -116 49 -82
<< metal1 >>
rect -9 -82 73 -72
rect -9 -116 15 -82
rect 49 -116 73 -82
rect -9 -126 73 -116
<< end >>
