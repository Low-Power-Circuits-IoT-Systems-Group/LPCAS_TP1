magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 75 151 80 200
rect 67 117 80 151
rect 75 83 80 117
rect 67 49 80 83
rect 75 0 80 49
<< nwell >>
rect -89 -36 111 362
<< pmos >>
rect 0 0 30 200
<< pdiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 151 75 200
rect 30 117 41 151
rect 30 83 75 117
rect 30 49 41 83
rect 30 0 75 49
<< pdiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
rect 41 117 75 151
rect 41 49 75 83
<< nsubdiff >>
rect -53 314 75 326
rect -53 280 -6 314
rect 28 280 75 314
rect -53 268 75 280
<< nsubdiffcont >>
rect -6 280 28 314
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -51 314 73 324
rect -51 280 -6 314
rect 28 280 73 314
rect -51 270 73 280
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
<< viali >>
rect -6 280 28 314
<< metal1 >>
rect -51 314 73 324
rect -51 280 -6 314
rect 28 280 73 314
rect -51 270 73 280
<< end >>
