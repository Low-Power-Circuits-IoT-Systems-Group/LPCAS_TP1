magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 1350
rect 611 0 650 1350
<< nwell >>
rect -47 -36 647 1512
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -11 0 0 1350
rect 600 0 611 1350
<< nsubdiff >>
rect -11 1464 611 1476
rect -11 1430 45 1464
rect 79 1430 113 1464
rect 147 1430 181 1464
rect 215 1430 249 1464
rect 283 1430 317 1464
rect 351 1430 385 1464
rect 419 1430 453 1464
rect 487 1430 521 1464
rect 555 1430 611 1464
rect -11 1418 611 1430
<< nsubdiffcont >>
rect 45 1430 79 1464
rect 113 1430 147 1464
rect 181 1430 215 1464
rect 249 1430 283 1464
rect 317 1430 351 1464
rect 385 1430 419 1464
rect 453 1430 487 1464
rect 521 1430 555 1464
<< poly >>
rect 0 1350 600 1380
rect 0 -30 600 0
<< locali >>
rect -9 1464 609 1474
rect -9 1430 31 1464
rect 79 1430 103 1464
rect 147 1430 175 1464
rect 215 1430 247 1464
rect 283 1430 317 1464
rect 353 1430 385 1464
rect 425 1430 453 1464
rect 497 1430 521 1464
rect 569 1430 609 1464
rect -9 1420 609 1430
<< viali >>
rect 31 1430 45 1464
rect 45 1430 65 1464
rect 103 1430 113 1464
rect 113 1430 137 1464
rect 175 1430 181 1464
rect 181 1430 209 1464
rect 247 1430 249 1464
rect 249 1430 281 1464
rect 319 1430 351 1464
rect 351 1430 353 1464
rect 391 1430 419 1464
rect 419 1430 425 1464
rect 463 1430 487 1464
rect 487 1430 497 1464
rect 535 1430 555 1464
rect 555 1430 569 1464
<< metal1 >>
rect -9 1464 609 1474
rect -9 1430 31 1464
rect 65 1430 103 1464
rect 137 1430 175 1464
rect 209 1430 247 1464
rect 281 1430 319 1464
rect 353 1430 391 1464
rect 425 1430 463 1464
rect 497 1430 535 1464
rect 569 1430 609 1464
rect -9 1420 609 1430
<< end >>
