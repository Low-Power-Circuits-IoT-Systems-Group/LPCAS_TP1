magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< pwell >>
rect -239 -26 1079 126
<< nmos >>
rect 0 0 1000 100
<< ndiff >>
rect -53 67 0 100
rect -53 33 -45 67
rect -11 33 0 67
rect -53 0 0 33
rect 1000 67 1053 100
rect 1000 33 1011 67
rect 1045 33 1053 67
rect 1000 0 1053 33
<< ndiffc >>
rect -45 33 -11 67
rect 1011 33 1045 67
<< psubdiff >>
rect -213 67 -107 100
rect -213 33 -177 67
rect -143 33 -107 67
rect -213 0 -107 33
<< psubdiffcont >>
rect -177 33 -143 67
<< poly >>
rect 0 182 1000 192
rect 0 148 16 182
rect 50 148 88 182
rect 122 148 160 182
rect 194 148 232 182
rect 266 148 304 182
rect 338 148 376 182
rect 410 148 448 182
rect 482 148 520 182
rect 554 148 592 182
rect 626 148 664 182
rect 698 148 736 182
rect 770 148 808 182
rect 842 148 879 182
rect 913 148 950 182
rect 984 148 1000 182
rect 0 100 1000 148
rect 0 -30 1000 0
<< polycont >>
rect 16 148 50 182
rect 88 148 122 182
rect 160 148 194 182
rect 232 148 266 182
rect 304 148 338 182
rect 376 148 410 182
rect 448 148 482 182
rect 520 148 554 182
rect 592 148 626 182
rect 664 148 698 182
rect 736 148 770 182
rect 808 148 842 182
rect 879 148 913 182
rect 950 148 984 182
<< locali >>
rect 0 182 1000 188
rect 0 148 16 182
rect 50 148 88 182
rect 128 148 160 182
rect 206 148 232 182
rect 284 148 304 182
rect 362 148 376 182
rect 440 148 448 182
rect 482 148 484 182
rect 518 148 520 182
rect 554 148 562 182
rect 626 148 640 182
rect 698 148 718 182
rect 770 148 796 182
rect 842 148 873 182
rect 913 148 950 182
rect 984 148 1000 182
rect 0 142 1000 148
rect -211 67 -109 100
rect -211 33 -177 67
rect -143 33 -109 67
rect -211 0 -109 33
rect -45 67 -11 100
rect -45 0 -11 33
rect 1011 67 1045 100
rect 1011 0 1045 33
<< viali >>
rect 16 148 50 182
rect 94 148 122 182
rect 122 148 128 182
rect 172 148 194 182
rect 194 148 206 182
rect 250 148 266 182
rect 266 148 284 182
rect 328 148 338 182
rect 338 148 362 182
rect 406 148 410 182
rect 410 148 440 182
rect 484 148 518 182
rect 562 148 592 182
rect 592 148 596 182
rect 640 148 664 182
rect 664 148 674 182
rect 718 148 736 182
rect 736 148 752 182
rect 796 148 808 182
rect 808 148 830 182
rect 873 148 879 182
rect 879 148 907 182
rect 950 148 984 182
rect -177 33 -143 67
<< metal1 >>
rect 0 182 1000 192
rect 0 148 16 182
rect 50 148 94 182
rect 128 148 172 182
rect 206 148 250 182
rect 284 148 328 182
rect 362 148 406 182
rect 440 148 484 182
rect 518 148 562 182
rect 596 148 640 182
rect 674 148 718 182
rect 752 148 796 182
rect 830 148 873 182
rect 907 148 950 182
rect 984 148 1000 182
rect 0 138 1000 148
rect -211 67 -109 100
rect -211 33 -177 67
rect -143 33 -109 67
rect -211 0 -109 33
<< end >>
