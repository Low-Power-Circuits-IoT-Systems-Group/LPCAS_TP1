magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< pwell >>
rect -79 -26 579 654
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -53 471 0 500
rect -53 437 -45 471
rect -11 437 0 471
rect -53 403 0 437
rect -53 369 -45 403
rect -11 369 0 403
rect -53 335 0 369
rect -53 301 -45 335
rect -11 301 0 335
rect -53 267 0 301
rect -53 233 -45 267
rect -11 233 0 267
rect -53 199 0 233
rect -53 165 -45 199
rect -11 165 0 199
rect -53 131 0 165
rect -53 97 -45 131
rect -11 97 0 131
rect -53 63 0 97
rect -53 29 -45 63
rect -11 29 0 63
rect -53 0 0 29
rect 500 471 553 500
rect 500 437 511 471
rect 545 437 553 471
rect 500 403 553 437
rect 500 369 511 403
rect 545 369 553 403
rect 500 335 553 369
rect 500 301 511 335
rect 545 301 553 335
rect 500 267 553 301
rect 500 233 511 267
rect 545 233 553 267
rect 500 199 553 233
rect 500 165 511 199
rect 545 165 553 199
rect 500 131 553 165
rect 500 97 511 131
rect 545 97 553 131
rect 500 63 553 97
rect 500 29 511 63
rect 545 29 553 63
rect 500 0 553 29
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< psubdiff >>
rect -53 616 553 628
rect -53 582 -5 616
rect 29 582 63 616
rect 97 582 131 616
rect 165 582 199 616
rect 233 582 267 616
rect 301 582 335 616
rect 369 582 403 616
rect 437 582 471 616
rect 505 582 553 616
rect -53 570 553 582
<< psubdiffcont >>
rect -5 582 29 616
rect 63 582 97 616
rect 131 582 165 616
rect 199 582 233 616
rect 267 582 301 616
rect 335 582 369 616
rect 403 582 437 616
rect 471 582 505 616
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect -51 616 551 626
rect -51 582 -19 616
rect 29 582 53 616
rect 97 582 125 616
rect 165 582 197 616
rect 233 582 267 616
rect 303 582 335 616
rect 375 582 403 616
rect 447 582 471 616
rect 519 582 551 616
rect -51 572 551 582
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
<< viali >>
rect -19 582 -5 616
rect -5 582 15 616
rect 53 582 63 616
rect 63 582 87 616
rect 125 582 131 616
rect 131 582 159 616
rect 197 582 199 616
rect 199 582 231 616
rect 269 582 301 616
rect 301 582 303 616
rect 341 582 369 616
rect 369 582 375 616
rect 413 582 437 616
rect 437 582 447 616
rect 485 582 505 616
rect 505 582 519 616
<< metal1 >>
rect -51 616 551 626
rect -51 582 -19 616
rect 15 582 53 616
rect 87 582 125 616
rect 159 582 197 616
rect 231 582 269 616
rect 303 582 341 616
rect 375 582 413 616
rect 447 582 485 616
rect 519 582 551 616
rect -51 572 551 582
<< end >>
