magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -64 26 64 27
rect -64 -26 -58 26
rect -6 -26 6 26
rect 58 -26 64 26
rect -64 -27 64 -26
<< via1 >>
rect -58 -26 -6 26
rect 6 -26 58 26
<< metal2 >>
rect -64 26 64 27
rect -64 -26 -58 26
rect -6 -26 6 26
rect 58 -26 64 26
rect -64 -27 64 -26
<< end >>
