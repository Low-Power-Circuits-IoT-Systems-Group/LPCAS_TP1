magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 471 -45 500
rect -50 437 -37 471
rect -50 403 -45 437
rect -50 369 -37 403
rect -50 335 -45 369
rect -50 301 -37 335
rect -50 267 -45 301
rect -50 233 -37 267
rect -50 199 -45 233
rect -50 165 -37 199
rect -50 131 -45 165
rect -50 97 -37 131
rect -50 63 -45 97
rect -50 29 -37 63
rect -50 0 -45 29
<< pwell >>
rect -71 -154 579 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -45 471 0 500
rect -11 437 0 471
rect -45 403 0 437
rect -11 369 0 403
rect -45 335 0 369
rect -11 301 0 335
rect -45 267 0 301
rect -11 233 0 267
rect -45 199 0 233
rect -11 165 0 199
rect -45 131 0 165
rect -11 97 0 131
rect -45 63 0 97
rect -11 29 0 63
rect -45 0 0 29
rect 500 471 553 500
rect 500 437 511 471
rect 545 437 553 471
rect 500 403 553 437
rect 500 369 511 403
rect 545 369 553 403
rect 500 335 553 369
rect 500 301 511 335
rect 545 301 553 335
rect 500 267 553 301
rect 500 233 511 267
rect 545 233 553 267
rect 500 199 553 233
rect 500 165 511 199
rect 545 165 553 199
rect 500 131 553 165
rect 500 97 511 131
rect 545 97 553 131
rect 500 63 553 97
rect 500 29 511 63
rect 545 29 553 63
rect 500 0 553 29
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< psubdiff >>
rect -45 -82 553 -70
rect -45 -116 -1 -82
rect 33 -116 67 -82
rect 101 -116 135 -82
rect 169 -116 203 -82
rect 237 -116 271 -82
rect 305 -116 339 -82
rect 373 -116 407 -82
rect 441 -116 475 -82
rect 509 -116 553 -82
rect -45 -128 553 -116
<< psubdiffcont >>
rect -1 -116 33 -82
rect 67 -116 101 -82
rect 135 -116 169 -82
rect 203 -116 237 -82
rect 271 -116 305 -82
rect 339 -116 373 -82
rect 407 -116 441 -82
rect 475 -116 509 -82
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
rect -43 -82 551 -72
rect -43 -116 -15 -82
rect 33 -116 57 -82
rect 101 -116 129 -82
rect 169 -116 201 -82
rect 237 -116 271 -82
rect 307 -116 339 -82
rect 379 -116 407 -82
rect 451 -116 475 -82
rect 523 -116 551 -82
rect -43 -126 551 -116
<< viali >>
rect -15 -116 -1 -82
rect -1 -116 19 -82
rect 57 -116 67 -82
rect 67 -116 91 -82
rect 129 -116 135 -82
rect 135 -116 163 -82
rect 201 -116 203 -82
rect 203 -116 235 -82
rect 273 -116 305 -82
rect 305 -116 307 -82
rect 345 -116 373 -82
rect 373 -116 379 -82
rect 417 -116 441 -82
rect 441 -116 451 -82
rect 489 -116 509 -82
rect 509 -116 523 -82
<< metal1 >>
rect -43 -82 551 -72
rect -43 -116 -15 -82
rect 19 -116 57 -82
rect 91 -116 129 -82
rect 163 -116 201 -82
rect 235 -116 273 -82
rect 307 -116 345 -82
rect 379 -116 417 -82
rect 451 -116 489 -82
rect 523 -116 551 -82
rect -43 -126 551 -116
<< end >>
