magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 0 0 19 1400
rect 311 0 330 1400
<< pwell >>
rect -37 -154 337 1426
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -11 0 0 1400
rect 300 0 311 1400
<< psubdiff >>
rect -11 -82 311 -70
rect -11 -116 31 -82
rect 65 -116 99 -82
rect 133 -116 167 -82
rect 201 -116 235 -82
rect 269 -116 311 -82
rect -11 -128 311 -116
<< psubdiffcont >>
rect 31 -116 65 -82
rect 99 -116 133 -82
rect 167 -116 201 -82
rect 235 -116 269 -82
<< poly >>
rect 0 1482 300 1492
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1400 300 1448
rect 0 -30 300 0
<< polycont >>
rect 16 1448 50 1482
rect 94 1448 128 1482
rect 172 1448 206 1482
rect 250 1448 284 1482
<< locali >>
rect 0 1482 300 1488
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1442 300 1448
rect -9 -82 309 -72
rect -9 -116 25 -82
rect 65 -116 97 -82
rect 133 -116 167 -82
rect 203 -116 235 -82
rect 275 -116 309 -82
rect -9 -126 309 -116
<< viali >>
rect 16 1448 50 1482
rect 94 1448 128 1482
rect 172 1448 206 1482
rect 250 1448 284 1482
rect 25 -116 31 -82
rect 31 -116 59 -82
rect 97 -116 99 -82
rect 99 -116 131 -82
rect 169 -116 201 -82
rect 201 -116 203 -82
rect 241 -116 269 -82
rect 269 -116 275 -82
<< metal1 >>
rect 0 1482 300 1492
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1438 300 1448
rect -9 -82 309 -72
rect -9 -116 25 -82
rect 59 -116 97 -82
rect 131 -116 169 -82
rect 203 -116 241 -82
rect 275 -116 309 -82
rect -9 -126 309 -116
<< end >>
