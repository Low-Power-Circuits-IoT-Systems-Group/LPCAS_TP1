magic
tech sky130A
timestamp 1741700111
<< metal1 >>
rect -13 61 13 64
rect -13 29 13 35
rect -13 -3 13 3
rect -13 -35 13 -29
rect -13 -64 13 -61
<< via1 >>
rect -13 35 13 61
rect -13 3 13 29
rect -13 -29 13 -3
rect -13 -61 13 -35
<< metal2 >>
rect -13 61 13 64
rect -13 29 13 35
rect -13 -3 13 3
rect -13 -35 13 -29
rect -13 -64 13 -61
<< end >>
