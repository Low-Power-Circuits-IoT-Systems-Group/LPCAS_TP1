magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< locali >>
rect -17 161 17 199
rect -17 89 17 127
rect -17 17 17 55
rect -17 -55 17 -17
rect -17 -127 17 -89
rect -17 -199 17 -161
<< viali >>
rect -17 199 17 233
rect -17 127 17 161
rect -17 55 17 89
rect -17 -17 17 17
rect -17 -89 17 -55
rect -17 -161 17 -127
rect -17 -233 17 -199
<< metal1 >>
rect -23 233 23 245
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -245 23 -233
<< end >>
