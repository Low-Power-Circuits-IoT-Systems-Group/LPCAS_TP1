magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 678 -45 710
rect -50 644 -37 678
rect -50 610 -45 644
rect -50 576 -37 610
rect -50 542 -45 576
rect -50 508 -37 542
rect -50 474 -45 508
rect -50 440 -37 474
rect -50 406 -45 440
rect -50 372 -37 406
rect -50 338 -45 372
rect -50 304 -37 338
rect -50 270 -45 304
rect -50 236 -37 270
rect -50 202 -45 236
rect -50 168 -37 202
rect -50 134 -45 168
rect -50 100 -37 134
rect -50 66 -45 100
rect -50 32 -37 66
rect -50 0 -45 32
<< nwell >>
rect -81 -36 289 872
<< pmos >>
rect 0 0 200 710
<< pdiff >>
rect -45 678 0 710
rect -11 644 0 678
rect -45 610 0 644
rect -11 576 0 610
rect -45 542 0 576
rect -11 508 0 542
rect -45 474 0 508
rect -11 440 0 474
rect -45 406 0 440
rect -11 372 0 406
rect -45 338 0 372
rect -11 304 0 338
rect -45 270 0 304
rect -11 236 0 270
rect -45 202 0 236
rect -11 168 0 202
rect -45 134 0 168
rect -11 100 0 134
rect -45 66 0 100
rect -11 32 0 66
rect -45 0 0 32
rect 200 678 253 710
rect 200 644 211 678
rect 245 644 253 678
rect 200 610 253 644
rect 200 576 211 610
rect 245 576 253 610
rect 200 542 253 576
rect 200 508 211 542
rect 245 508 253 542
rect 200 474 253 508
rect 200 440 211 474
rect 245 440 253 474
rect 200 406 253 440
rect 200 372 211 406
rect 245 372 253 406
rect 200 338 253 372
rect 200 304 211 338
rect 245 304 253 338
rect 200 270 253 304
rect 200 236 211 270
rect 245 236 253 270
rect 200 202 253 236
rect 200 168 211 202
rect 245 168 253 202
rect 200 134 253 168
rect 200 100 211 134
rect 245 100 253 134
rect 200 66 253 100
rect 200 32 211 66
rect 245 32 253 66
rect 200 0 253 32
<< pdiffc >>
rect -45 644 -11 678
rect -45 576 -11 610
rect -45 508 -11 542
rect -45 440 -11 474
rect -45 372 -11 406
rect -45 304 -11 338
rect -45 236 -11 270
rect -45 168 -11 202
rect -45 100 -11 134
rect -45 32 -11 66
rect 211 644 245 678
rect 211 576 245 610
rect 211 508 245 542
rect 211 440 245 474
rect 211 372 245 406
rect 211 304 245 338
rect 211 236 245 270
rect 211 168 245 202
rect 211 100 245 134
rect 211 32 245 66
<< nsubdiff >>
rect -45 824 253 836
rect -45 790 -15 824
rect 19 790 53 824
rect 87 790 121 824
rect 155 790 189 824
rect 223 790 253 824
rect -45 778 253 790
<< nsubdiffcont >>
rect -15 790 19 824
rect 53 790 87 824
rect 121 790 155 824
rect 189 790 223 824
<< poly >>
rect 0 710 200 740
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect -43 824 251 834
rect -43 790 -21 824
rect 19 790 51 824
rect 87 790 121 824
rect 157 790 189 824
rect 229 790 251 824
rect -43 780 251 790
rect -45 678 -11 710
rect -45 610 -11 644
rect -45 542 -11 576
rect -45 474 -11 508
rect -45 406 -11 440
rect -45 338 -11 372
rect -45 270 -11 304
rect -45 202 -11 236
rect -45 134 -11 168
rect -45 66 -11 100
rect -45 0 -11 32
rect 211 678 245 710
rect 211 610 245 644
rect 211 542 245 576
rect 211 474 245 508
rect 211 406 245 440
rect 211 338 245 372
rect 211 270 245 304
rect 211 202 245 236
rect 211 134 245 168
rect 211 66 245 100
rect 211 0 245 32
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect -21 790 -15 824
rect -15 790 13 824
rect 51 790 53 824
rect 53 790 85 824
rect 123 790 155 824
rect 155 790 157 824
rect 195 790 223 824
rect 223 790 229 824
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect -43 824 251 834
rect -43 790 -21 824
rect 13 790 51 824
rect 85 790 123 824
rect 157 790 195 824
rect 229 790 251 824
rect -43 780 251 790
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
