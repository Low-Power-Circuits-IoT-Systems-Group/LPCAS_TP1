magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< pwell >>
rect -79 -154 109 226
<< nmos >>
rect 0 0 30 200
<< ndiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 151 83 200
rect 30 117 41 151
rect 75 117 83 151
rect 30 83 83 117
rect 30 49 41 83
rect 75 49 83 83
rect 30 0 83 49
<< ndiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
rect 41 117 75 151
rect 41 49 75 83
<< psubdiff >>
rect -53 -82 83 -70
rect -53 -116 -2 -82
rect 32 -116 83 -82
rect -53 -128 83 -116
<< psubdiffcont >>
rect -2 -116 32 -82
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
rect -51 -82 81 -72
rect -51 -116 -2 -82
rect 32 -116 81 -82
rect -51 -126 81 -116
<< viali >>
rect -2 -116 32 -82
<< metal1 >>
rect -51 -82 81 -72
rect -51 -116 -2 -82
rect 32 -116 81 -82
rect -51 -126 81 -116
<< end >>
