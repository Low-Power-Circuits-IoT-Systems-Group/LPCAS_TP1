magic
tech sky130A
timestamp 1741700111
<< metal1 >>
rect -13 125 13 128
rect -13 93 13 99
rect -13 61 13 67
rect -13 29 13 35
rect -13 -3 13 3
rect -13 -35 13 -29
rect -13 -67 13 -61
rect -13 -99 13 -93
rect -13 -128 13 -125
<< via1 >>
rect -13 99 13 125
rect -13 67 13 93
rect -13 35 13 61
rect -13 3 13 29
rect -13 -29 13 -3
rect -13 -61 13 -35
rect -13 -93 13 -67
rect -13 -125 13 -99
<< metal2 >>
rect -13 125 13 128
rect -13 93 13 99
rect -13 61 13 67
rect -13 29 13 35
rect -13 -3 13 3
rect -13 -35 13 -29
rect -13 -67 13 -61
rect -13 -99 13 -93
rect -13 -128 13 -125
<< end >>
