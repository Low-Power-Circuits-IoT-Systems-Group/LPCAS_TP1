magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 41 0 80 200
<< pwell >>
rect -79 -154 67 226
<< nmos >>
rect 0 0 30 200
<< ndiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 0 41 200
<< ndiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
<< psubdiff >>
rect -53 -82 41 -70
rect -53 -116 -23 -82
rect 11 -116 41 -82
rect -53 -128 41 -116
<< psubdiffcont >>
rect -23 -116 11 -82
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
rect -51 -82 39 -72
rect -51 -116 -23 -82
rect 11 -116 39 -82
rect -51 -126 39 -116
<< viali >>
rect -23 -116 11 -82
<< metal1 >>
rect -51 -82 39 -72
rect -51 -116 -23 -82
rect 11 -116 39 -82
rect -51 -126 39 -116
<< end >>
