magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -37 -32 -26 20
rect 26 -32 37 20
<< via1 >>
rect -26 -32 26 20
<< metal2 >>
rect -50 -32 -26 20
rect 26 -32 50 20
<< end >>
