magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< nwell >>
rect -89 -36 689 837
<< pmos >>
rect 0 0 600 675
<< pdiff >>
rect -53 626 0 675
rect -53 592 -45 626
rect -11 592 0 626
rect -53 558 0 592
rect -53 524 -45 558
rect -11 524 0 558
rect -53 490 0 524
rect -53 456 -45 490
rect -11 456 0 490
rect -53 422 0 456
rect -53 388 -45 422
rect -11 388 0 422
rect -53 354 0 388
rect -53 320 -45 354
rect -11 320 0 354
rect -53 286 0 320
rect -53 252 -45 286
rect -11 252 0 286
rect -53 218 0 252
rect -53 184 -45 218
rect -11 184 0 218
rect -53 150 0 184
rect -53 116 -45 150
rect -11 116 0 150
rect -53 82 0 116
rect -53 48 -45 82
rect -11 48 0 82
rect -53 0 0 48
rect 600 626 653 675
rect 600 592 611 626
rect 645 592 653 626
rect 600 558 653 592
rect 600 524 611 558
rect 645 524 653 558
rect 600 490 653 524
rect 600 456 611 490
rect 645 456 653 490
rect 600 422 653 456
rect 600 388 611 422
rect 645 388 653 422
rect 600 354 653 388
rect 600 320 611 354
rect 645 320 653 354
rect 600 286 653 320
rect 600 252 611 286
rect 645 252 653 286
rect 600 218 653 252
rect 600 184 611 218
rect 645 184 653 218
rect 600 150 653 184
rect 600 116 611 150
rect 645 116 653 150
rect 600 82 653 116
rect 600 48 611 82
rect 645 48 653 82
rect 600 0 653 48
<< pdiffc >>
rect -45 592 -11 626
rect -45 524 -11 558
rect -45 456 -11 490
rect -45 388 -11 422
rect -45 320 -11 354
rect -45 252 -11 286
rect -45 184 -11 218
rect -45 116 -11 150
rect -45 48 -11 82
rect 611 592 645 626
rect 611 524 645 558
rect 611 456 645 490
rect 611 388 645 422
rect 611 320 645 354
rect 611 252 645 286
rect 611 184 645 218
rect 611 116 645 150
rect 611 48 645 82
<< nsubdiff >>
rect -53 789 653 801
rect -53 755 -23 789
rect 11 755 45 789
rect 79 755 113 789
rect 147 755 181 789
rect 215 755 249 789
rect 283 755 317 789
rect 351 755 385 789
rect 419 755 453 789
rect 487 755 521 789
rect 555 755 589 789
rect 623 755 653 789
rect -53 743 653 755
<< nsubdiffcont >>
rect -23 755 11 789
rect 45 755 79 789
rect 113 755 147 789
rect 181 755 215 789
rect 249 755 283 789
rect 317 755 351 789
rect 385 755 419 789
rect 453 755 487 789
rect 521 755 555 789
rect 589 755 623 789
<< poly >>
rect 0 675 600 705
rect 0 -48 600 0
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< polycont >>
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< locali >>
rect -51 789 651 799
rect -51 755 -23 789
rect 29 755 45 789
rect 101 755 113 789
rect 173 755 181 789
rect 245 755 249 789
rect 351 755 355 789
rect 419 755 427 789
rect 487 755 499 789
rect 555 755 571 789
rect 623 755 651 789
rect -51 745 651 755
rect -45 626 -11 675
rect -45 558 -11 592
rect -45 490 -11 524
rect -45 422 -11 456
rect -45 354 -11 388
rect -45 286 -11 320
rect -45 218 -11 252
rect -45 150 -11 184
rect -45 82 -11 116
rect -45 0 -11 48
rect 611 626 645 675
rect 611 558 645 592
rect 611 490 645 524
rect 611 422 645 456
rect 611 354 645 388
rect 611 286 645 320
rect 611 218 645 252
rect 611 150 645 184
rect 611 82 645 116
rect 611 0 645 48
rect 0 -48 600 -42
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -88 600 -82
<< viali >>
rect -5 755 11 789
rect 11 755 29 789
rect 67 755 79 789
rect 79 755 101 789
rect 139 755 147 789
rect 147 755 173 789
rect 211 755 215 789
rect 215 755 245 789
rect 283 755 317 789
rect 355 755 385 789
rect 385 755 389 789
rect 427 755 453 789
rect 453 755 461 789
rect 499 755 521 789
rect 521 755 533 789
rect 571 755 589 789
rect 589 755 605 789
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< metal1 >>
rect -51 789 651 799
rect -51 755 -5 789
rect 29 755 67 789
rect 101 755 139 789
rect 173 755 211 789
rect 245 755 283 789
rect 317 755 355 789
rect 389 755 427 789
rect 461 755 499 789
rect 533 755 571 789
rect 605 755 651 789
rect -51 745 651 755
rect 0 -48 600 -38
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< end >>
