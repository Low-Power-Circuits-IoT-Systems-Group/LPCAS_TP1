magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 1350
rect 645 1304 650 1350
rect 637 1270 650 1304
rect 645 1236 650 1270
rect 637 1202 650 1236
rect 645 1168 650 1202
rect 637 1134 650 1168
rect 645 1100 650 1134
rect 637 1066 650 1100
rect 645 1032 650 1066
rect 637 998 650 1032
rect 645 964 650 998
rect 637 930 650 964
rect 645 896 650 930
rect 637 862 650 896
rect 645 828 650 862
rect 637 794 650 828
rect 645 760 650 794
rect 637 726 650 760
rect 645 692 650 726
rect 637 658 650 692
rect 645 624 650 658
rect 637 590 650 624
rect 645 556 650 590
rect 637 522 650 556
rect 645 488 650 522
rect 637 454 650 488
rect 645 420 650 454
rect 637 386 650 420
rect 645 352 650 386
rect 637 318 650 352
rect 645 284 650 318
rect 637 250 650 284
rect 645 216 650 250
rect 637 182 650 216
rect 645 148 650 182
rect 637 114 650 148
rect 645 80 650 114
rect 637 46 650 80
rect 645 0 650 46
<< nwell >>
rect -47 -36 681 1512
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -11 0 0 1350
rect 600 1304 645 1350
rect 600 1270 611 1304
rect 600 1236 645 1270
rect 600 1202 611 1236
rect 600 1168 645 1202
rect 600 1134 611 1168
rect 600 1100 645 1134
rect 600 1066 611 1100
rect 600 1032 645 1066
rect 600 998 611 1032
rect 600 964 645 998
rect 600 930 611 964
rect 600 896 645 930
rect 600 862 611 896
rect 600 828 645 862
rect 600 794 611 828
rect 600 760 645 794
rect 600 726 611 760
rect 600 692 645 726
rect 600 658 611 692
rect 600 624 645 658
rect 600 590 611 624
rect 600 556 645 590
rect 600 522 611 556
rect 600 488 645 522
rect 600 454 611 488
rect 600 420 645 454
rect 600 386 611 420
rect 600 352 645 386
rect 600 318 611 352
rect 600 284 645 318
rect 600 250 611 284
rect 600 216 645 250
rect 600 182 611 216
rect 600 148 645 182
rect 600 114 611 148
rect 600 80 645 114
rect 600 46 611 80
rect 600 0 645 46
<< pdiffc >>
rect 611 1270 645 1304
rect 611 1202 645 1236
rect 611 1134 645 1168
rect 611 1066 645 1100
rect 611 998 645 1032
rect 611 930 645 964
rect 611 862 645 896
rect 611 794 645 828
rect 611 726 645 760
rect 611 658 645 692
rect 611 590 645 624
rect 611 522 645 556
rect 611 454 645 488
rect 611 386 645 420
rect 611 318 645 352
rect 611 250 645 284
rect 611 182 645 216
rect 611 114 645 148
rect 611 46 645 80
<< nsubdiff >>
rect -11 1464 645 1476
rect -11 1430 28 1464
rect 62 1430 96 1464
rect 130 1430 164 1464
rect 198 1430 232 1464
rect 266 1430 300 1464
rect 334 1430 368 1464
rect 402 1430 436 1464
rect 470 1430 504 1464
rect 538 1430 572 1464
rect 606 1430 645 1464
rect -11 1418 645 1430
<< nsubdiffcont >>
rect 28 1430 62 1464
rect 96 1430 130 1464
rect 164 1430 198 1464
rect 232 1430 266 1464
rect 300 1430 334 1464
rect 368 1430 402 1464
rect 436 1430 470 1464
rect 504 1430 538 1464
rect 572 1430 606 1464
<< poly >>
rect 0 1350 600 1380
rect 0 -30 600 0
<< locali >>
rect -9 1464 643 1474
rect -9 1430 12 1464
rect 62 1430 84 1464
rect 130 1430 156 1464
rect 198 1430 228 1464
rect 266 1430 300 1464
rect 334 1430 368 1464
rect 406 1430 436 1464
rect 478 1430 504 1464
rect 550 1430 572 1464
rect 622 1430 643 1464
rect -9 1420 643 1430
rect 611 1304 645 1350
rect 611 1236 645 1270
rect 611 1168 645 1202
rect 611 1100 645 1134
rect 611 1032 645 1066
rect 611 964 645 998
rect 611 896 645 930
rect 611 828 645 862
rect 611 760 645 794
rect 611 692 645 726
rect 611 624 645 658
rect 611 556 645 590
rect 611 488 645 522
rect 611 420 645 454
rect 611 352 645 386
rect 611 284 645 318
rect 611 216 645 250
rect 611 148 645 182
rect 611 80 645 114
rect 611 0 645 46
<< viali >>
rect 12 1430 28 1464
rect 28 1430 46 1464
rect 84 1430 96 1464
rect 96 1430 118 1464
rect 156 1430 164 1464
rect 164 1430 190 1464
rect 228 1430 232 1464
rect 232 1430 262 1464
rect 300 1430 334 1464
rect 372 1430 402 1464
rect 402 1430 406 1464
rect 444 1430 470 1464
rect 470 1430 478 1464
rect 516 1430 538 1464
rect 538 1430 550 1464
rect 588 1430 606 1464
rect 606 1430 622 1464
<< metal1 >>
rect -9 1464 643 1474
rect -9 1430 12 1464
rect 46 1430 84 1464
rect 118 1430 156 1464
rect 190 1430 228 1464
rect 262 1430 300 1464
rect 334 1430 372 1464
rect 406 1430 444 1464
rect 478 1430 516 1464
rect 550 1430 588 1464
rect 622 1430 643 1464
rect -9 1420 643 1430
<< end >>
