magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< nwell >>
rect -89 -36 689 1512
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -53 1304 0 1350
rect -53 1270 -45 1304
rect -11 1270 0 1304
rect -53 1236 0 1270
rect -53 1202 -45 1236
rect -11 1202 0 1236
rect -53 1168 0 1202
rect -53 1134 -45 1168
rect -11 1134 0 1168
rect -53 1100 0 1134
rect -53 1066 -45 1100
rect -11 1066 0 1100
rect -53 1032 0 1066
rect -53 998 -45 1032
rect -11 998 0 1032
rect -53 964 0 998
rect -53 930 -45 964
rect -11 930 0 964
rect -53 896 0 930
rect -53 862 -45 896
rect -11 862 0 896
rect -53 828 0 862
rect -53 794 -45 828
rect -11 794 0 828
rect -53 760 0 794
rect -53 726 -45 760
rect -11 726 0 760
rect -53 692 0 726
rect -53 658 -45 692
rect -11 658 0 692
rect -53 624 0 658
rect -53 590 -45 624
rect -11 590 0 624
rect -53 556 0 590
rect -53 522 -45 556
rect -11 522 0 556
rect -53 488 0 522
rect -53 454 -45 488
rect -11 454 0 488
rect -53 420 0 454
rect -53 386 -45 420
rect -11 386 0 420
rect -53 352 0 386
rect -53 318 -45 352
rect -11 318 0 352
rect -53 284 0 318
rect -53 250 -45 284
rect -11 250 0 284
rect -53 216 0 250
rect -53 182 -45 216
rect -11 182 0 216
rect -53 148 0 182
rect -53 114 -45 148
rect -11 114 0 148
rect -53 80 0 114
rect -53 46 -45 80
rect -11 46 0 80
rect -53 0 0 46
rect 600 1304 653 1350
rect 600 1270 611 1304
rect 645 1270 653 1304
rect 600 1236 653 1270
rect 600 1202 611 1236
rect 645 1202 653 1236
rect 600 1168 653 1202
rect 600 1134 611 1168
rect 645 1134 653 1168
rect 600 1100 653 1134
rect 600 1066 611 1100
rect 645 1066 653 1100
rect 600 1032 653 1066
rect 600 998 611 1032
rect 645 998 653 1032
rect 600 964 653 998
rect 600 930 611 964
rect 645 930 653 964
rect 600 896 653 930
rect 600 862 611 896
rect 645 862 653 896
rect 600 828 653 862
rect 600 794 611 828
rect 645 794 653 828
rect 600 760 653 794
rect 600 726 611 760
rect 645 726 653 760
rect 600 692 653 726
rect 600 658 611 692
rect 645 658 653 692
rect 600 624 653 658
rect 600 590 611 624
rect 645 590 653 624
rect 600 556 653 590
rect 600 522 611 556
rect 645 522 653 556
rect 600 488 653 522
rect 600 454 611 488
rect 645 454 653 488
rect 600 420 653 454
rect 600 386 611 420
rect 645 386 653 420
rect 600 352 653 386
rect 600 318 611 352
rect 645 318 653 352
rect 600 284 653 318
rect 600 250 611 284
rect 645 250 653 284
rect 600 216 653 250
rect 600 182 611 216
rect 645 182 653 216
rect 600 148 653 182
rect 600 114 611 148
rect 645 114 653 148
rect 600 80 653 114
rect 600 46 611 80
rect 645 46 653 80
rect 600 0 653 46
<< pdiffc >>
rect -45 1270 -11 1304
rect -45 1202 -11 1236
rect -45 1134 -11 1168
rect -45 1066 -11 1100
rect -45 998 -11 1032
rect -45 930 -11 964
rect -45 862 -11 896
rect -45 794 -11 828
rect -45 726 -11 760
rect -45 658 -11 692
rect -45 590 -11 624
rect -45 522 -11 556
rect -45 454 -11 488
rect -45 386 -11 420
rect -45 318 -11 352
rect -45 250 -11 284
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect 611 1270 645 1304
rect 611 1202 645 1236
rect 611 1134 645 1168
rect 611 1066 645 1100
rect 611 998 645 1032
rect 611 930 645 964
rect 611 862 645 896
rect 611 794 645 828
rect 611 726 645 760
rect 611 658 645 692
rect 611 590 645 624
rect 611 522 645 556
rect 611 454 645 488
rect 611 386 645 420
rect 611 318 645 352
rect 611 250 645 284
rect 611 182 645 216
rect 611 114 645 148
rect 611 46 645 80
<< nsubdiff >>
rect -53 1464 653 1476
rect -53 1430 -23 1464
rect 11 1430 45 1464
rect 79 1430 113 1464
rect 147 1430 181 1464
rect 215 1430 249 1464
rect 283 1430 317 1464
rect 351 1430 385 1464
rect 419 1430 453 1464
rect 487 1430 521 1464
rect 555 1430 589 1464
rect 623 1430 653 1464
rect -53 1418 653 1430
<< nsubdiffcont >>
rect -23 1430 11 1464
rect 45 1430 79 1464
rect 113 1430 147 1464
rect 181 1430 215 1464
rect 249 1430 283 1464
rect 317 1430 351 1464
rect 385 1430 419 1464
rect 453 1430 487 1464
rect 521 1430 555 1464
rect 589 1430 623 1464
<< poly >>
rect 0 1350 600 1380
rect 0 -30 600 0
<< locali >>
rect -51 1464 651 1474
rect -51 1430 -23 1464
rect 29 1430 45 1464
rect 101 1430 113 1464
rect 173 1430 181 1464
rect 245 1430 249 1464
rect 351 1430 355 1464
rect 419 1430 427 1464
rect 487 1430 499 1464
rect 555 1430 571 1464
rect 623 1430 651 1464
rect -51 1420 651 1430
rect -45 1304 -11 1350
rect -45 1236 -11 1270
rect -45 1168 -11 1202
rect -45 1100 -11 1134
rect -45 1032 -11 1066
rect -45 964 -11 998
rect -45 896 -11 930
rect -45 828 -11 862
rect -45 760 -11 794
rect -45 692 -11 726
rect -45 624 -11 658
rect -45 556 -11 590
rect -45 488 -11 522
rect -45 420 -11 454
rect -45 352 -11 386
rect -45 284 -11 318
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 0 -11 46
rect 611 1304 645 1350
rect 611 1236 645 1270
rect 611 1168 645 1202
rect 611 1100 645 1134
rect 611 1032 645 1066
rect 611 964 645 998
rect 611 896 645 930
rect 611 828 645 862
rect 611 760 645 794
rect 611 692 645 726
rect 611 624 645 658
rect 611 556 645 590
rect 611 488 645 522
rect 611 420 645 454
rect 611 352 645 386
rect 611 284 645 318
rect 611 216 645 250
rect 611 148 645 182
rect 611 80 645 114
rect 611 0 645 46
<< viali >>
rect -5 1430 11 1464
rect 11 1430 29 1464
rect 67 1430 79 1464
rect 79 1430 101 1464
rect 139 1430 147 1464
rect 147 1430 173 1464
rect 211 1430 215 1464
rect 215 1430 245 1464
rect 283 1430 317 1464
rect 355 1430 385 1464
rect 385 1430 389 1464
rect 427 1430 453 1464
rect 453 1430 461 1464
rect 499 1430 521 1464
rect 521 1430 533 1464
rect 571 1430 589 1464
rect 589 1430 605 1464
<< metal1 >>
rect -51 1464 651 1474
rect -51 1430 -5 1464
rect 29 1430 67 1464
rect 101 1430 139 1464
rect 173 1430 211 1464
rect 245 1430 283 1464
rect 317 1430 355 1464
rect 389 1430 427 1464
rect 461 1430 499 1464
rect 533 1430 571 1464
rect 605 1430 651 1464
rect -51 1420 651 1430
<< end >>
