magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -17 -17 17 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -55 17 55 23
rect -55 -17 -17 17
rect 17 -17 55 17
rect -55 -23 55 -17
<< end >>
