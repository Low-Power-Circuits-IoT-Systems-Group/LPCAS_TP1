magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -17 -17 17 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -26 17 26 32
rect -26 -17 -17 17
rect 17 -17 26 17
rect -26 -32 26 -17
<< end >>
