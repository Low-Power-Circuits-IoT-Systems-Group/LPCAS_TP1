magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< locali >>
rect -17 269 17 307
rect -17 197 17 235
rect -17 125 17 163
rect -17 53 17 91
rect -17 -19 17 19
rect -17 -91 17 -53
rect -17 -163 17 -125
rect -17 -235 17 -197
rect -17 -307 17 -269
<< viali >>
rect -17 307 17 341
rect -17 235 17 269
rect -17 163 17 197
rect -17 91 17 125
rect -17 19 17 53
rect -17 -53 17 -19
rect -17 -125 17 -91
rect -17 -197 17 -163
rect -17 -269 17 -235
rect -17 -341 17 -307
<< metal1 >>
rect -23 341 23 353
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -353 23 -341
<< end >>
