magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< xpolycontact >>
rect -141 253 141 685
rect -141 -685 141 -253
<< xpolyres >>
rect -141 -253 141 253
<< viali >>
rect -125 271 125 665
rect -125 -666 125 -272
<< metal1 >>
rect -131 665 131 679
rect -131 271 -125 665
rect 125 271 131 665
rect -131 258 131 271
rect -131 -272 131 -258
rect -131 -666 -125 -272
rect 125 -666 131 -272
rect -131 -679 131 -666
<< end >>
