magic
tech sky130A
magscale 1 2
timestamp 1748330293
<< nwell >>
rect 6916 33585 7962 34758
rect 9409 34388 23891 37672
rect 6916 33187 8118 33585
rect 6916 33185 7962 33187
rect 9409 33164 16229 34388
rect 8928 15209 9974 16382
rect 11421 16012 25903 19296
rect 8928 14811 10130 15209
rect 8928 14809 9974 14811
rect 11421 14788 18241 16012
<< pwell >>
rect 7612 33118 7950 33124
rect 6926 33066 8062 33118
rect 6926 33032 8098 33066
rect 6926 31958 7012 33032
rect 7976 32980 8098 33032
rect 6828 31872 7012 31958
rect 6828 31625 6914 31872
rect 6828 31539 7420 31625
rect 7334 30994 7420 31539
rect 7305 30908 7420 30994
rect 8012 30994 8098 32980
rect 9408 32978 16402 33064
rect 9408 31612 14404 32978
rect 16316 31612 16402 32978
rect 9408 31526 16402 31612
rect 9408 31368 11302 31526
rect 9408 31106 9494 31368
rect 11216 31106 11302 31368
rect 8012 30908 8127 30994
rect 7305 30709 7391 30908
rect 8041 30709 8127 30908
rect 7305 30623 8127 30709
rect 9408 29410 11302 31106
rect 12642 31320 14646 31526
rect 12642 31110 12728 31320
rect 14560 31110 14646 31320
rect 12642 31024 14646 31110
rect 9624 14742 9962 14748
rect 8938 14690 10074 14742
rect 8938 14656 10110 14690
rect 8938 13582 9024 14656
rect 9988 14604 10110 14656
rect 8840 13496 9024 13582
rect 8840 13249 8926 13496
rect 8840 13163 9432 13249
rect 9346 12618 9432 13163
rect 9317 12532 9432 12618
rect 10024 12618 10110 14604
rect 11420 14602 18414 14688
rect 10024 12532 10139 12618
rect 9317 12333 9403 12532
rect 10053 12333 10139 12532
rect 9317 12247 10139 12333
rect 11420 11120 11506 14602
rect 13228 13236 13402 14602
rect 18328 13236 18414 14602
rect 13228 13150 18414 13236
rect 13228 11120 13314 13150
rect 11420 11034 13314 11120
<< nmos >>
rect 11495 32348 11995 32848
rect 12051 32348 12551 32848
rect 12607 32348 13107 32848
rect 13269 32348 13769 32848
rect 13825 32348 14325 32848
rect 11495 31794 11995 32294
rect 12051 31794 12551 32294
rect 12607 31794 13107 32294
rect 13269 31794 13769 32294
rect 13825 31794 14325 32294
<< pmos >>
rect 9622 36036 10222 37386
rect 10384 36036 10984 37386
rect 11040 36036 11640 37386
rect 11696 36036 12296 37386
rect 12352 36036 12952 37386
rect 13008 36036 13608 37386
rect 13664 36036 14264 37386
rect 9622 34614 10222 35964
rect 10384 34614 10984 35964
rect 11040 34614 11640 35964
rect 11696 34614 12296 35964
rect 12352 34614 12952 35964
rect 13008 34614 13608 35964
rect 13664 34614 14264 35964
rect 19132 36018 19732 37368
rect 19788 36018 20388 37368
rect 20444 36018 21044 37368
rect 21100 36018 21700 37368
rect 21756 36018 22356 37368
rect 22412 36018 23012 37368
rect 9820 33499 10020 34099
rect 10076 33499 10276 34099
rect 10332 33499 10532 34099
rect 10694 33499 10894 34099
rect 10950 33499 11150 34099
rect 11206 33499 11406 34099
rect 12008 33414 12208 34124
rect 12264 33414 12464 34124
rect 12520 33414 12720 34124
rect 13142 33431 13742 34106
rect 13920 33431 14520 34106
<< nmoslvt >>
rect 9674 31394 9974 32794
rect 10030 31394 10330 32794
rect 10386 31394 10686 32794
rect 10742 31394 11042 32794
rect 9674 29680 9974 31080
rect 10030 29680 10330 31080
rect 10386 29680 10686 31080
rect 10742 29680 11042 31080
<< ndiff >>
rect 9621 32757 9674 32794
rect 9621 32723 9629 32757
rect 9663 32723 9674 32757
rect 9621 32689 9674 32723
rect 9621 32655 9629 32689
rect 9663 32655 9674 32689
rect 9621 32621 9674 32655
rect 9621 32587 9629 32621
rect 9663 32587 9674 32621
rect 9621 32553 9674 32587
rect 9621 32519 9629 32553
rect 9663 32519 9674 32553
rect 9621 32485 9674 32519
rect 9621 32451 9629 32485
rect 9663 32451 9674 32485
rect 9621 32417 9674 32451
rect 9621 32383 9629 32417
rect 9663 32383 9674 32417
rect 9621 32349 9674 32383
rect 9621 32315 9629 32349
rect 9663 32315 9674 32349
rect 9621 32281 9674 32315
rect 9621 32247 9629 32281
rect 9663 32247 9674 32281
rect 9621 32213 9674 32247
rect 9621 32179 9629 32213
rect 9663 32179 9674 32213
rect 9621 32145 9674 32179
rect 9621 32111 9629 32145
rect 9663 32111 9674 32145
rect 9621 32077 9674 32111
rect 9621 32043 9629 32077
rect 9663 32043 9674 32077
rect 9621 32009 9674 32043
rect 9621 31975 9629 32009
rect 9663 31975 9674 32009
rect 9621 31941 9674 31975
rect 9621 31907 9629 31941
rect 9663 31907 9674 31941
rect 9621 31873 9674 31907
rect 9621 31839 9629 31873
rect 9663 31839 9674 31873
rect 9621 31805 9674 31839
rect 9621 31771 9629 31805
rect 9663 31771 9674 31805
rect 9621 31737 9674 31771
rect 9621 31703 9629 31737
rect 9663 31703 9674 31737
rect 9621 31669 9674 31703
rect 9621 31635 9629 31669
rect 9663 31635 9674 31669
rect 9621 31601 9674 31635
rect 9621 31567 9629 31601
rect 9663 31567 9674 31601
rect 9621 31533 9674 31567
rect 9621 31499 9629 31533
rect 9663 31499 9674 31533
rect 9621 31465 9674 31499
rect 9621 31431 9629 31465
rect 9663 31431 9674 31465
rect 9621 31394 9674 31431
rect 9974 32757 10030 32794
rect 9974 32723 9985 32757
rect 10019 32723 10030 32757
rect 9974 32689 10030 32723
rect 9974 32655 9985 32689
rect 10019 32655 10030 32689
rect 9974 32621 10030 32655
rect 9974 32587 9985 32621
rect 10019 32587 10030 32621
rect 9974 32553 10030 32587
rect 9974 32519 9985 32553
rect 10019 32519 10030 32553
rect 9974 32485 10030 32519
rect 9974 32451 9985 32485
rect 10019 32451 10030 32485
rect 9974 32417 10030 32451
rect 9974 32383 9985 32417
rect 10019 32383 10030 32417
rect 9974 32349 10030 32383
rect 9974 32315 9985 32349
rect 10019 32315 10030 32349
rect 9974 32281 10030 32315
rect 9974 32247 9985 32281
rect 10019 32247 10030 32281
rect 9974 32213 10030 32247
rect 9974 32179 9985 32213
rect 10019 32179 10030 32213
rect 9974 32145 10030 32179
rect 9974 32111 9985 32145
rect 10019 32111 10030 32145
rect 9974 32077 10030 32111
rect 9974 32043 9985 32077
rect 10019 32043 10030 32077
rect 9974 32009 10030 32043
rect 9974 31975 9985 32009
rect 10019 31975 10030 32009
rect 9974 31941 10030 31975
rect 9974 31907 9985 31941
rect 10019 31907 10030 31941
rect 9974 31873 10030 31907
rect 9974 31839 9985 31873
rect 10019 31839 10030 31873
rect 9974 31805 10030 31839
rect 9974 31771 9985 31805
rect 10019 31771 10030 31805
rect 9974 31737 10030 31771
rect 9974 31703 9985 31737
rect 10019 31703 10030 31737
rect 9974 31669 10030 31703
rect 9974 31635 9985 31669
rect 10019 31635 10030 31669
rect 9974 31601 10030 31635
rect 9974 31567 9985 31601
rect 10019 31567 10030 31601
rect 9974 31533 10030 31567
rect 9974 31499 9985 31533
rect 10019 31499 10030 31533
rect 9974 31465 10030 31499
rect 9974 31431 9985 31465
rect 10019 31431 10030 31465
rect 9974 31394 10030 31431
rect 10330 32757 10386 32794
rect 10330 32723 10341 32757
rect 10375 32723 10386 32757
rect 10330 32689 10386 32723
rect 10330 32655 10341 32689
rect 10375 32655 10386 32689
rect 10330 32621 10386 32655
rect 10330 32587 10341 32621
rect 10375 32587 10386 32621
rect 10330 32553 10386 32587
rect 10330 32519 10341 32553
rect 10375 32519 10386 32553
rect 10330 32485 10386 32519
rect 10330 32451 10341 32485
rect 10375 32451 10386 32485
rect 10330 32417 10386 32451
rect 10330 32383 10341 32417
rect 10375 32383 10386 32417
rect 10330 32349 10386 32383
rect 10330 32315 10341 32349
rect 10375 32315 10386 32349
rect 10330 32281 10386 32315
rect 10330 32247 10341 32281
rect 10375 32247 10386 32281
rect 10330 32213 10386 32247
rect 10330 32179 10341 32213
rect 10375 32179 10386 32213
rect 10330 32145 10386 32179
rect 10330 32111 10341 32145
rect 10375 32111 10386 32145
rect 10330 32077 10386 32111
rect 10330 32043 10341 32077
rect 10375 32043 10386 32077
rect 10330 32009 10386 32043
rect 10330 31975 10341 32009
rect 10375 31975 10386 32009
rect 10330 31941 10386 31975
rect 10330 31907 10341 31941
rect 10375 31907 10386 31941
rect 10330 31873 10386 31907
rect 10330 31839 10341 31873
rect 10375 31839 10386 31873
rect 10330 31805 10386 31839
rect 10330 31771 10341 31805
rect 10375 31771 10386 31805
rect 10330 31737 10386 31771
rect 10330 31703 10341 31737
rect 10375 31703 10386 31737
rect 10330 31669 10386 31703
rect 10330 31635 10341 31669
rect 10375 31635 10386 31669
rect 10330 31601 10386 31635
rect 10330 31567 10341 31601
rect 10375 31567 10386 31601
rect 10330 31533 10386 31567
rect 10330 31499 10341 31533
rect 10375 31499 10386 31533
rect 10330 31465 10386 31499
rect 10330 31431 10341 31465
rect 10375 31431 10386 31465
rect 10330 31394 10386 31431
rect 10686 32757 10742 32794
rect 10686 32723 10697 32757
rect 10731 32723 10742 32757
rect 10686 32689 10742 32723
rect 10686 32655 10697 32689
rect 10731 32655 10742 32689
rect 10686 32621 10742 32655
rect 10686 32587 10697 32621
rect 10731 32587 10742 32621
rect 10686 32553 10742 32587
rect 10686 32519 10697 32553
rect 10731 32519 10742 32553
rect 10686 32485 10742 32519
rect 10686 32451 10697 32485
rect 10731 32451 10742 32485
rect 10686 32417 10742 32451
rect 10686 32383 10697 32417
rect 10731 32383 10742 32417
rect 10686 32349 10742 32383
rect 10686 32315 10697 32349
rect 10731 32315 10742 32349
rect 10686 32281 10742 32315
rect 10686 32247 10697 32281
rect 10731 32247 10742 32281
rect 10686 32213 10742 32247
rect 10686 32179 10697 32213
rect 10731 32179 10742 32213
rect 10686 32145 10742 32179
rect 10686 32111 10697 32145
rect 10731 32111 10742 32145
rect 10686 32077 10742 32111
rect 10686 32043 10697 32077
rect 10731 32043 10742 32077
rect 10686 32009 10742 32043
rect 10686 31975 10697 32009
rect 10731 31975 10742 32009
rect 10686 31941 10742 31975
rect 10686 31907 10697 31941
rect 10731 31907 10742 31941
rect 10686 31873 10742 31907
rect 10686 31839 10697 31873
rect 10731 31839 10742 31873
rect 10686 31805 10742 31839
rect 10686 31771 10697 31805
rect 10731 31771 10742 31805
rect 10686 31737 10742 31771
rect 10686 31703 10697 31737
rect 10731 31703 10742 31737
rect 10686 31669 10742 31703
rect 10686 31635 10697 31669
rect 10731 31635 10742 31669
rect 10686 31601 10742 31635
rect 10686 31567 10697 31601
rect 10731 31567 10742 31601
rect 10686 31533 10742 31567
rect 10686 31499 10697 31533
rect 10731 31499 10742 31533
rect 10686 31465 10742 31499
rect 10686 31431 10697 31465
rect 10731 31431 10742 31465
rect 10686 31394 10742 31431
rect 11042 32757 11095 32794
rect 11042 32723 11053 32757
rect 11087 32723 11095 32757
rect 11042 32689 11095 32723
rect 11042 32655 11053 32689
rect 11087 32655 11095 32689
rect 11042 32621 11095 32655
rect 11042 32587 11053 32621
rect 11087 32587 11095 32621
rect 11042 32553 11095 32587
rect 11042 32519 11053 32553
rect 11087 32519 11095 32553
rect 11042 32485 11095 32519
rect 11042 32451 11053 32485
rect 11087 32451 11095 32485
rect 11042 32417 11095 32451
rect 11042 32383 11053 32417
rect 11087 32383 11095 32417
rect 11042 32349 11095 32383
rect 11042 32315 11053 32349
rect 11087 32315 11095 32349
rect 11042 32281 11095 32315
rect 11042 32247 11053 32281
rect 11087 32247 11095 32281
rect 11042 32213 11095 32247
rect 11042 32179 11053 32213
rect 11087 32179 11095 32213
rect 11042 32145 11095 32179
rect 11042 32111 11053 32145
rect 11087 32111 11095 32145
rect 11042 32077 11095 32111
rect 11042 32043 11053 32077
rect 11087 32043 11095 32077
rect 11042 32009 11095 32043
rect 11042 31975 11053 32009
rect 11087 31975 11095 32009
rect 11042 31941 11095 31975
rect 11042 31907 11053 31941
rect 11087 31907 11095 31941
rect 11042 31873 11095 31907
rect 11042 31839 11053 31873
rect 11087 31839 11095 31873
rect 11042 31805 11095 31839
rect 11042 31771 11053 31805
rect 11087 31771 11095 31805
rect 11042 31737 11095 31771
rect 11042 31703 11053 31737
rect 11087 31703 11095 31737
rect 11042 31669 11095 31703
rect 11042 31635 11053 31669
rect 11087 31635 11095 31669
rect 11042 31601 11095 31635
rect 11042 31567 11053 31601
rect 11087 31567 11095 31601
rect 11042 31533 11095 31567
rect 11042 31499 11053 31533
rect 11087 31499 11095 31533
rect 11042 31465 11095 31499
rect 11042 31431 11053 31465
rect 11087 31431 11095 31465
rect 11042 31394 11095 31431
rect 11442 32819 11495 32848
rect 11442 32785 11450 32819
rect 11484 32785 11495 32819
rect 11442 32751 11495 32785
rect 11442 32717 11450 32751
rect 11484 32717 11495 32751
rect 11442 32683 11495 32717
rect 11442 32649 11450 32683
rect 11484 32649 11495 32683
rect 11442 32615 11495 32649
rect 11442 32581 11450 32615
rect 11484 32581 11495 32615
rect 11442 32547 11495 32581
rect 11442 32513 11450 32547
rect 11484 32513 11495 32547
rect 11442 32479 11495 32513
rect 11442 32445 11450 32479
rect 11484 32445 11495 32479
rect 11442 32411 11495 32445
rect 11442 32377 11450 32411
rect 11484 32377 11495 32411
rect 11442 32348 11495 32377
rect 11995 32819 12051 32848
rect 11995 32785 12006 32819
rect 12040 32785 12051 32819
rect 11995 32751 12051 32785
rect 11995 32717 12006 32751
rect 12040 32717 12051 32751
rect 11995 32683 12051 32717
rect 11995 32649 12006 32683
rect 12040 32649 12051 32683
rect 11995 32615 12051 32649
rect 11995 32581 12006 32615
rect 12040 32581 12051 32615
rect 11995 32547 12051 32581
rect 11995 32513 12006 32547
rect 12040 32513 12051 32547
rect 11995 32479 12051 32513
rect 11995 32445 12006 32479
rect 12040 32445 12051 32479
rect 11995 32411 12051 32445
rect 11995 32377 12006 32411
rect 12040 32377 12051 32411
rect 11995 32348 12051 32377
rect 12551 32819 12607 32848
rect 12551 32785 12562 32819
rect 12596 32785 12607 32819
rect 12551 32751 12607 32785
rect 12551 32717 12562 32751
rect 12596 32717 12607 32751
rect 12551 32683 12607 32717
rect 12551 32649 12562 32683
rect 12596 32649 12607 32683
rect 12551 32615 12607 32649
rect 12551 32581 12562 32615
rect 12596 32581 12607 32615
rect 12551 32547 12607 32581
rect 12551 32513 12562 32547
rect 12596 32513 12607 32547
rect 12551 32479 12607 32513
rect 12551 32445 12562 32479
rect 12596 32445 12607 32479
rect 12551 32411 12607 32445
rect 12551 32377 12562 32411
rect 12596 32377 12607 32411
rect 12551 32348 12607 32377
rect 13107 32819 13160 32848
rect 13107 32785 13118 32819
rect 13152 32785 13160 32819
rect 13107 32751 13160 32785
rect 13107 32717 13118 32751
rect 13152 32717 13160 32751
rect 13107 32683 13160 32717
rect 13107 32649 13118 32683
rect 13152 32649 13160 32683
rect 13107 32615 13160 32649
rect 13107 32581 13118 32615
rect 13152 32581 13160 32615
rect 13107 32547 13160 32581
rect 13107 32513 13118 32547
rect 13152 32513 13160 32547
rect 13107 32479 13160 32513
rect 13107 32445 13118 32479
rect 13152 32445 13160 32479
rect 13107 32411 13160 32445
rect 13107 32377 13118 32411
rect 13152 32377 13160 32411
rect 13107 32348 13160 32377
rect 13216 32819 13269 32848
rect 13216 32785 13224 32819
rect 13258 32785 13269 32819
rect 13216 32751 13269 32785
rect 13216 32717 13224 32751
rect 13258 32717 13269 32751
rect 13216 32683 13269 32717
rect 13216 32649 13224 32683
rect 13258 32649 13269 32683
rect 13216 32615 13269 32649
rect 13216 32581 13224 32615
rect 13258 32581 13269 32615
rect 13216 32547 13269 32581
rect 13216 32513 13224 32547
rect 13258 32513 13269 32547
rect 13216 32479 13269 32513
rect 13216 32445 13224 32479
rect 13258 32445 13269 32479
rect 13216 32411 13269 32445
rect 13216 32377 13224 32411
rect 13258 32377 13269 32411
rect 13216 32348 13269 32377
rect 13769 32819 13825 32848
rect 13769 32785 13780 32819
rect 13814 32785 13825 32819
rect 13769 32751 13825 32785
rect 13769 32717 13780 32751
rect 13814 32717 13825 32751
rect 13769 32683 13825 32717
rect 13769 32649 13780 32683
rect 13814 32649 13825 32683
rect 13769 32615 13825 32649
rect 13769 32581 13780 32615
rect 13814 32581 13825 32615
rect 13769 32547 13825 32581
rect 13769 32513 13780 32547
rect 13814 32513 13825 32547
rect 13769 32479 13825 32513
rect 13769 32445 13780 32479
rect 13814 32445 13825 32479
rect 13769 32411 13825 32445
rect 13769 32377 13780 32411
rect 13814 32377 13825 32411
rect 13769 32348 13825 32377
rect 14325 32819 14378 32848
rect 14325 32785 14336 32819
rect 14370 32785 14378 32819
rect 14325 32751 14378 32785
rect 14325 32717 14336 32751
rect 14370 32717 14378 32751
rect 14325 32683 14378 32717
rect 14325 32649 14336 32683
rect 14370 32649 14378 32683
rect 14325 32615 14378 32649
rect 14325 32581 14336 32615
rect 14370 32581 14378 32615
rect 14325 32547 14378 32581
rect 14325 32513 14336 32547
rect 14370 32513 14378 32547
rect 14325 32479 14378 32513
rect 14325 32445 14336 32479
rect 14370 32445 14378 32479
rect 14325 32411 14378 32445
rect 14325 32377 14336 32411
rect 14370 32377 14378 32411
rect 14325 32348 14378 32377
rect 11442 32265 11495 32294
rect 11442 32231 11450 32265
rect 11484 32231 11495 32265
rect 11442 32197 11495 32231
rect 11442 32163 11450 32197
rect 11484 32163 11495 32197
rect 11442 32129 11495 32163
rect 11442 32095 11450 32129
rect 11484 32095 11495 32129
rect 11442 32061 11495 32095
rect 11442 32027 11450 32061
rect 11484 32027 11495 32061
rect 11442 31993 11495 32027
rect 11442 31959 11450 31993
rect 11484 31959 11495 31993
rect 11442 31925 11495 31959
rect 11442 31891 11450 31925
rect 11484 31891 11495 31925
rect 11442 31857 11495 31891
rect 11442 31823 11450 31857
rect 11484 31823 11495 31857
rect 11442 31794 11495 31823
rect 11995 32265 12051 32294
rect 11995 32231 12006 32265
rect 12040 32231 12051 32265
rect 11995 32197 12051 32231
rect 11995 32163 12006 32197
rect 12040 32163 12051 32197
rect 11995 32129 12051 32163
rect 11995 32095 12006 32129
rect 12040 32095 12051 32129
rect 11995 32061 12051 32095
rect 11995 32027 12006 32061
rect 12040 32027 12051 32061
rect 11995 31993 12051 32027
rect 11995 31959 12006 31993
rect 12040 31959 12051 31993
rect 11995 31925 12051 31959
rect 11995 31891 12006 31925
rect 12040 31891 12051 31925
rect 11995 31857 12051 31891
rect 11995 31823 12006 31857
rect 12040 31823 12051 31857
rect 11995 31794 12051 31823
rect 12551 32265 12607 32294
rect 12551 32231 12562 32265
rect 12596 32231 12607 32265
rect 12551 32197 12607 32231
rect 12551 32163 12562 32197
rect 12596 32163 12607 32197
rect 12551 32129 12607 32163
rect 12551 32095 12562 32129
rect 12596 32095 12607 32129
rect 12551 32061 12607 32095
rect 12551 32027 12562 32061
rect 12596 32027 12607 32061
rect 12551 31993 12607 32027
rect 12551 31959 12562 31993
rect 12596 31959 12607 31993
rect 12551 31925 12607 31959
rect 12551 31891 12562 31925
rect 12596 31891 12607 31925
rect 12551 31857 12607 31891
rect 12551 31823 12562 31857
rect 12596 31823 12607 31857
rect 12551 31794 12607 31823
rect 13107 32265 13160 32294
rect 13107 32231 13118 32265
rect 13152 32231 13160 32265
rect 13107 32197 13160 32231
rect 13107 32163 13118 32197
rect 13152 32163 13160 32197
rect 13107 32129 13160 32163
rect 13107 32095 13118 32129
rect 13152 32095 13160 32129
rect 13107 32061 13160 32095
rect 13107 32027 13118 32061
rect 13152 32027 13160 32061
rect 13107 31993 13160 32027
rect 13107 31959 13118 31993
rect 13152 31959 13160 31993
rect 13107 31925 13160 31959
rect 13107 31891 13118 31925
rect 13152 31891 13160 31925
rect 13107 31857 13160 31891
rect 13107 31823 13118 31857
rect 13152 31823 13160 31857
rect 13107 31794 13160 31823
rect 13216 32265 13269 32294
rect 13216 32231 13224 32265
rect 13258 32231 13269 32265
rect 13216 32197 13269 32231
rect 13216 32163 13224 32197
rect 13258 32163 13269 32197
rect 13216 32129 13269 32163
rect 13216 32095 13224 32129
rect 13258 32095 13269 32129
rect 13216 32061 13269 32095
rect 13216 32027 13224 32061
rect 13258 32027 13269 32061
rect 13216 31993 13269 32027
rect 13216 31959 13224 31993
rect 13258 31959 13269 31993
rect 13216 31925 13269 31959
rect 13216 31891 13224 31925
rect 13258 31891 13269 31925
rect 13216 31857 13269 31891
rect 13216 31823 13224 31857
rect 13258 31823 13269 31857
rect 13216 31794 13269 31823
rect 13769 32265 13825 32294
rect 13769 32231 13780 32265
rect 13814 32231 13825 32265
rect 13769 32197 13825 32231
rect 13769 32163 13780 32197
rect 13814 32163 13825 32197
rect 13769 32129 13825 32163
rect 13769 32095 13780 32129
rect 13814 32095 13825 32129
rect 13769 32061 13825 32095
rect 13769 32027 13780 32061
rect 13814 32027 13825 32061
rect 13769 31993 13825 32027
rect 13769 31959 13780 31993
rect 13814 31959 13825 31993
rect 13769 31925 13825 31959
rect 13769 31891 13780 31925
rect 13814 31891 13825 31925
rect 13769 31857 13825 31891
rect 13769 31823 13780 31857
rect 13814 31823 13825 31857
rect 13769 31794 13825 31823
rect 14325 32265 14378 32294
rect 14325 32231 14336 32265
rect 14370 32231 14378 32265
rect 14325 32197 14378 32231
rect 14325 32163 14336 32197
rect 14370 32163 14378 32197
rect 14325 32129 14378 32163
rect 14325 32095 14336 32129
rect 14370 32095 14378 32129
rect 14325 32061 14378 32095
rect 14325 32027 14336 32061
rect 14370 32027 14378 32061
rect 14325 31993 14378 32027
rect 14325 31959 14336 31993
rect 14370 31959 14378 31993
rect 14325 31925 14378 31959
rect 14325 31891 14336 31925
rect 14370 31891 14378 31925
rect 14325 31857 14378 31891
rect 14325 31823 14336 31857
rect 14370 31823 14378 31857
rect 14325 31794 14378 31823
rect 9621 31043 9674 31080
rect 9621 31009 9629 31043
rect 9663 31009 9674 31043
rect 9621 30975 9674 31009
rect 9621 30941 9629 30975
rect 9663 30941 9674 30975
rect 9621 30907 9674 30941
rect 9621 30873 9629 30907
rect 9663 30873 9674 30907
rect 9621 30839 9674 30873
rect 9621 30805 9629 30839
rect 9663 30805 9674 30839
rect 9621 30771 9674 30805
rect 9621 30737 9629 30771
rect 9663 30737 9674 30771
rect 9621 30703 9674 30737
rect 9621 30669 9629 30703
rect 9663 30669 9674 30703
rect 9621 30635 9674 30669
rect 9621 30601 9629 30635
rect 9663 30601 9674 30635
rect 9621 30567 9674 30601
rect 9621 30533 9629 30567
rect 9663 30533 9674 30567
rect 9621 30499 9674 30533
rect 9621 30465 9629 30499
rect 9663 30465 9674 30499
rect 9621 30431 9674 30465
rect 9621 30397 9629 30431
rect 9663 30397 9674 30431
rect 9621 30363 9674 30397
rect 9621 30329 9629 30363
rect 9663 30329 9674 30363
rect 9621 30295 9674 30329
rect 9621 30261 9629 30295
rect 9663 30261 9674 30295
rect 9621 30227 9674 30261
rect 9621 30193 9629 30227
rect 9663 30193 9674 30227
rect 9621 30159 9674 30193
rect 9621 30125 9629 30159
rect 9663 30125 9674 30159
rect 9621 30091 9674 30125
rect 9621 30057 9629 30091
rect 9663 30057 9674 30091
rect 9621 30023 9674 30057
rect 9621 29989 9629 30023
rect 9663 29989 9674 30023
rect 9621 29955 9674 29989
rect 9621 29921 9629 29955
rect 9663 29921 9674 29955
rect 9621 29887 9674 29921
rect 9621 29853 9629 29887
rect 9663 29853 9674 29887
rect 9621 29819 9674 29853
rect 9621 29785 9629 29819
rect 9663 29785 9674 29819
rect 9621 29751 9674 29785
rect 9621 29717 9629 29751
rect 9663 29717 9674 29751
rect 9621 29680 9674 29717
rect 9974 31043 10030 31080
rect 9974 31009 9985 31043
rect 10019 31009 10030 31043
rect 9974 30975 10030 31009
rect 9974 30941 9985 30975
rect 10019 30941 10030 30975
rect 9974 30907 10030 30941
rect 9974 30873 9985 30907
rect 10019 30873 10030 30907
rect 9974 30839 10030 30873
rect 9974 30805 9985 30839
rect 10019 30805 10030 30839
rect 9974 30771 10030 30805
rect 9974 30737 9985 30771
rect 10019 30737 10030 30771
rect 9974 30703 10030 30737
rect 9974 30669 9985 30703
rect 10019 30669 10030 30703
rect 9974 30635 10030 30669
rect 9974 30601 9985 30635
rect 10019 30601 10030 30635
rect 9974 30567 10030 30601
rect 9974 30533 9985 30567
rect 10019 30533 10030 30567
rect 9974 30499 10030 30533
rect 9974 30465 9985 30499
rect 10019 30465 10030 30499
rect 9974 30431 10030 30465
rect 9974 30397 9985 30431
rect 10019 30397 10030 30431
rect 9974 30363 10030 30397
rect 9974 30329 9985 30363
rect 10019 30329 10030 30363
rect 9974 30295 10030 30329
rect 9974 30261 9985 30295
rect 10019 30261 10030 30295
rect 9974 30227 10030 30261
rect 9974 30193 9985 30227
rect 10019 30193 10030 30227
rect 9974 30159 10030 30193
rect 9974 30125 9985 30159
rect 10019 30125 10030 30159
rect 9974 30091 10030 30125
rect 9974 30057 9985 30091
rect 10019 30057 10030 30091
rect 9974 30023 10030 30057
rect 9974 29989 9985 30023
rect 10019 29989 10030 30023
rect 9974 29955 10030 29989
rect 9974 29921 9985 29955
rect 10019 29921 10030 29955
rect 9974 29887 10030 29921
rect 9974 29853 9985 29887
rect 10019 29853 10030 29887
rect 9974 29819 10030 29853
rect 9974 29785 9985 29819
rect 10019 29785 10030 29819
rect 9974 29751 10030 29785
rect 9974 29717 9985 29751
rect 10019 29717 10030 29751
rect 9974 29680 10030 29717
rect 10330 31043 10386 31080
rect 10330 31009 10341 31043
rect 10375 31009 10386 31043
rect 10330 30975 10386 31009
rect 10330 30941 10341 30975
rect 10375 30941 10386 30975
rect 10330 30907 10386 30941
rect 10330 30873 10341 30907
rect 10375 30873 10386 30907
rect 10330 30839 10386 30873
rect 10330 30805 10341 30839
rect 10375 30805 10386 30839
rect 10330 30771 10386 30805
rect 10330 30737 10341 30771
rect 10375 30737 10386 30771
rect 10330 30703 10386 30737
rect 10330 30669 10341 30703
rect 10375 30669 10386 30703
rect 10330 30635 10386 30669
rect 10330 30601 10341 30635
rect 10375 30601 10386 30635
rect 10330 30567 10386 30601
rect 10330 30533 10341 30567
rect 10375 30533 10386 30567
rect 10330 30499 10386 30533
rect 10330 30465 10341 30499
rect 10375 30465 10386 30499
rect 10330 30431 10386 30465
rect 10330 30397 10341 30431
rect 10375 30397 10386 30431
rect 10330 30363 10386 30397
rect 10330 30329 10341 30363
rect 10375 30329 10386 30363
rect 10330 30295 10386 30329
rect 10330 30261 10341 30295
rect 10375 30261 10386 30295
rect 10330 30227 10386 30261
rect 10330 30193 10341 30227
rect 10375 30193 10386 30227
rect 10330 30159 10386 30193
rect 10330 30125 10341 30159
rect 10375 30125 10386 30159
rect 10330 30091 10386 30125
rect 10330 30057 10341 30091
rect 10375 30057 10386 30091
rect 10330 30023 10386 30057
rect 10330 29989 10341 30023
rect 10375 29989 10386 30023
rect 10330 29955 10386 29989
rect 10330 29921 10341 29955
rect 10375 29921 10386 29955
rect 10330 29887 10386 29921
rect 10330 29853 10341 29887
rect 10375 29853 10386 29887
rect 10330 29819 10386 29853
rect 10330 29785 10341 29819
rect 10375 29785 10386 29819
rect 10330 29751 10386 29785
rect 10330 29717 10341 29751
rect 10375 29717 10386 29751
rect 10330 29680 10386 29717
rect 10686 31043 10742 31080
rect 10686 31009 10697 31043
rect 10731 31009 10742 31043
rect 10686 30975 10742 31009
rect 10686 30941 10697 30975
rect 10731 30941 10742 30975
rect 10686 30907 10742 30941
rect 10686 30873 10697 30907
rect 10731 30873 10742 30907
rect 10686 30839 10742 30873
rect 10686 30805 10697 30839
rect 10731 30805 10742 30839
rect 10686 30771 10742 30805
rect 10686 30737 10697 30771
rect 10731 30737 10742 30771
rect 10686 30703 10742 30737
rect 10686 30669 10697 30703
rect 10731 30669 10742 30703
rect 10686 30635 10742 30669
rect 10686 30601 10697 30635
rect 10731 30601 10742 30635
rect 10686 30567 10742 30601
rect 10686 30533 10697 30567
rect 10731 30533 10742 30567
rect 10686 30499 10742 30533
rect 10686 30465 10697 30499
rect 10731 30465 10742 30499
rect 10686 30431 10742 30465
rect 10686 30397 10697 30431
rect 10731 30397 10742 30431
rect 10686 30363 10742 30397
rect 10686 30329 10697 30363
rect 10731 30329 10742 30363
rect 10686 30295 10742 30329
rect 10686 30261 10697 30295
rect 10731 30261 10742 30295
rect 10686 30227 10742 30261
rect 10686 30193 10697 30227
rect 10731 30193 10742 30227
rect 10686 30159 10742 30193
rect 10686 30125 10697 30159
rect 10731 30125 10742 30159
rect 10686 30091 10742 30125
rect 10686 30057 10697 30091
rect 10731 30057 10742 30091
rect 10686 30023 10742 30057
rect 10686 29989 10697 30023
rect 10731 29989 10742 30023
rect 10686 29955 10742 29989
rect 10686 29921 10697 29955
rect 10731 29921 10742 29955
rect 10686 29887 10742 29921
rect 10686 29853 10697 29887
rect 10731 29853 10742 29887
rect 10686 29819 10742 29853
rect 10686 29785 10697 29819
rect 10731 29785 10742 29819
rect 10686 29751 10742 29785
rect 10686 29717 10697 29751
rect 10731 29717 10742 29751
rect 10686 29680 10742 29717
rect 11042 31043 11095 31080
rect 11042 31009 11053 31043
rect 11087 31009 11095 31043
rect 11042 30975 11095 31009
rect 11042 30941 11053 30975
rect 11087 30941 11095 30975
rect 11042 30907 11095 30941
rect 11042 30873 11053 30907
rect 11087 30873 11095 30907
rect 11042 30839 11095 30873
rect 11042 30805 11053 30839
rect 11087 30805 11095 30839
rect 11042 30771 11095 30805
rect 11042 30737 11053 30771
rect 11087 30737 11095 30771
rect 11042 30703 11095 30737
rect 11042 30669 11053 30703
rect 11087 30669 11095 30703
rect 11042 30635 11095 30669
rect 11042 30601 11053 30635
rect 11087 30601 11095 30635
rect 11042 30567 11095 30601
rect 11042 30533 11053 30567
rect 11087 30533 11095 30567
rect 11042 30499 11095 30533
rect 11042 30465 11053 30499
rect 11087 30465 11095 30499
rect 11042 30431 11095 30465
rect 11042 30397 11053 30431
rect 11087 30397 11095 30431
rect 11042 30363 11095 30397
rect 11042 30329 11053 30363
rect 11087 30329 11095 30363
rect 11042 30295 11095 30329
rect 11042 30261 11053 30295
rect 11087 30261 11095 30295
rect 11042 30227 11095 30261
rect 11042 30193 11053 30227
rect 11087 30193 11095 30227
rect 11042 30159 11095 30193
rect 11042 30125 11053 30159
rect 11087 30125 11095 30159
rect 11042 30091 11095 30125
rect 11042 30057 11053 30091
rect 11087 30057 11095 30091
rect 11042 30023 11095 30057
rect 11042 29989 11053 30023
rect 11087 29989 11095 30023
rect 11042 29955 11095 29989
rect 11042 29921 11053 29955
rect 11087 29921 11095 29955
rect 11042 29887 11095 29921
rect 11042 29853 11053 29887
rect 11087 29853 11095 29887
rect 11042 29819 11095 29853
rect 11042 29785 11053 29819
rect 11087 29785 11095 29819
rect 11042 29751 11095 29785
rect 11042 29717 11053 29751
rect 11087 29717 11095 29751
rect 11042 29680 11095 29717
<< pdiff >>
rect 9569 37340 9622 37386
rect 9569 37306 9577 37340
rect 9611 37306 9622 37340
rect 9569 37272 9622 37306
rect 9569 37238 9577 37272
rect 9611 37238 9622 37272
rect 9569 37204 9622 37238
rect 9569 37170 9577 37204
rect 9611 37170 9622 37204
rect 9569 37136 9622 37170
rect 9569 37102 9577 37136
rect 9611 37102 9622 37136
rect 9569 37068 9622 37102
rect 9569 37034 9577 37068
rect 9611 37034 9622 37068
rect 9569 37000 9622 37034
rect 9569 36966 9577 37000
rect 9611 36966 9622 37000
rect 9569 36932 9622 36966
rect 9569 36898 9577 36932
rect 9611 36898 9622 36932
rect 9569 36864 9622 36898
rect 9569 36830 9577 36864
rect 9611 36830 9622 36864
rect 9569 36796 9622 36830
rect 9569 36762 9577 36796
rect 9611 36762 9622 36796
rect 9569 36728 9622 36762
rect 9569 36694 9577 36728
rect 9611 36694 9622 36728
rect 9569 36660 9622 36694
rect 9569 36626 9577 36660
rect 9611 36626 9622 36660
rect 9569 36592 9622 36626
rect 9569 36558 9577 36592
rect 9611 36558 9622 36592
rect 9569 36524 9622 36558
rect 9569 36490 9577 36524
rect 9611 36490 9622 36524
rect 9569 36456 9622 36490
rect 9569 36422 9577 36456
rect 9611 36422 9622 36456
rect 9569 36388 9622 36422
rect 9569 36354 9577 36388
rect 9611 36354 9622 36388
rect 9569 36320 9622 36354
rect 9569 36286 9577 36320
rect 9611 36286 9622 36320
rect 9569 36252 9622 36286
rect 9569 36218 9577 36252
rect 9611 36218 9622 36252
rect 9569 36184 9622 36218
rect 9569 36150 9577 36184
rect 9611 36150 9622 36184
rect 9569 36116 9622 36150
rect 9569 36082 9577 36116
rect 9611 36082 9622 36116
rect 9569 36036 9622 36082
rect 10222 37340 10275 37386
rect 10222 37306 10233 37340
rect 10267 37306 10275 37340
rect 10222 37272 10275 37306
rect 10222 37238 10233 37272
rect 10267 37238 10275 37272
rect 10222 37204 10275 37238
rect 10222 37170 10233 37204
rect 10267 37170 10275 37204
rect 10222 37136 10275 37170
rect 10222 37102 10233 37136
rect 10267 37102 10275 37136
rect 10222 37068 10275 37102
rect 10222 37034 10233 37068
rect 10267 37034 10275 37068
rect 10222 37000 10275 37034
rect 10222 36966 10233 37000
rect 10267 36966 10275 37000
rect 10222 36932 10275 36966
rect 10222 36898 10233 36932
rect 10267 36898 10275 36932
rect 10222 36864 10275 36898
rect 10222 36830 10233 36864
rect 10267 36830 10275 36864
rect 10222 36796 10275 36830
rect 10222 36762 10233 36796
rect 10267 36762 10275 36796
rect 10222 36728 10275 36762
rect 10222 36694 10233 36728
rect 10267 36694 10275 36728
rect 10222 36660 10275 36694
rect 10222 36626 10233 36660
rect 10267 36626 10275 36660
rect 10222 36592 10275 36626
rect 10222 36558 10233 36592
rect 10267 36558 10275 36592
rect 10222 36524 10275 36558
rect 10222 36490 10233 36524
rect 10267 36490 10275 36524
rect 10222 36456 10275 36490
rect 10222 36422 10233 36456
rect 10267 36422 10275 36456
rect 10222 36388 10275 36422
rect 10222 36354 10233 36388
rect 10267 36354 10275 36388
rect 10222 36320 10275 36354
rect 10222 36286 10233 36320
rect 10267 36286 10275 36320
rect 10222 36252 10275 36286
rect 10222 36218 10233 36252
rect 10267 36218 10275 36252
rect 10222 36184 10275 36218
rect 10222 36150 10233 36184
rect 10267 36150 10275 36184
rect 10222 36116 10275 36150
rect 10222 36082 10233 36116
rect 10267 36082 10275 36116
rect 10222 36036 10275 36082
rect 10331 37340 10384 37386
rect 10331 37306 10339 37340
rect 10373 37306 10384 37340
rect 10331 37272 10384 37306
rect 10331 37238 10339 37272
rect 10373 37238 10384 37272
rect 10331 37204 10384 37238
rect 10331 37170 10339 37204
rect 10373 37170 10384 37204
rect 10331 37136 10384 37170
rect 10331 37102 10339 37136
rect 10373 37102 10384 37136
rect 10331 37068 10384 37102
rect 10331 37034 10339 37068
rect 10373 37034 10384 37068
rect 10331 37000 10384 37034
rect 10331 36966 10339 37000
rect 10373 36966 10384 37000
rect 10331 36932 10384 36966
rect 10331 36898 10339 36932
rect 10373 36898 10384 36932
rect 10331 36864 10384 36898
rect 10331 36830 10339 36864
rect 10373 36830 10384 36864
rect 10331 36796 10384 36830
rect 10331 36762 10339 36796
rect 10373 36762 10384 36796
rect 10331 36728 10384 36762
rect 10331 36694 10339 36728
rect 10373 36694 10384 36728
rect 10331 36660 10384 36694
rect 10331 36626 10339 36660
rect 10373 36626 10384 36660
rect 10331 36592 10384 36626
rect 10331 36558 10339 36592
rect 10373 36558 10384 36592
rect 10331 36524 10384 36558
rect 10331 36490 10339 36524
rect 10373 36490 10384 36524
rect 10331 36456 10384 36490
rect 10331 36422 10339 36456
rect 10373 36422 10384 36456
rect 10331 36388 10384 36422
rect 10331 36354 10339 36388
rect 10373 36354 10384 36388
rect 10331 36320 10384 36354
rect 10331 36286 10339 36320
rect 10373 36286 10384 36320
rect 10331 36252 10384 36286
rect 10331 36218 10339 36252
rect 10373 36218 10384 36252
rect 10331 36184 10384 36218
rect 10331 36150 10339 36184
rect 10373 36150 10384 36184
rect 10331 36116 10384 36150
rect 10331 36082 10339 36116
rect 10373 36082 10384 36116
rect 10331 36036 10384 36082
rect 10984 37340 11040 37386
rect 10984 37306 10995 37340
rect 11029 37306 11040 37340
rect 10984 37272 11040 37306
rect 10984 37238 10995 37272
rect 11029 37238 11040 37272
rect 10984 37204 11040 37238
rect 10984 37170 10995 37204
rect 11029 37170 11040 37204
rect 10984 37136 11040 37170
rect 10984 37102 10995 37136
rect 11029 37102 11040 37136
rect 10984 37068 11040 37102
rect 10984 37034 10995 37068
rect 11029 37034 11040 37068
rect 10984 37000 11040 37034
rect 10984 36966 10995 37000
rect 11029 36966 11040 37000
rect 10984 36932 11040 36966
rect 10984 36898 10995 36932
rect 11029 36898 11040 36932
rect 10984 36864 11040 36898
rect 10984 36830 10995 36864
rect 11029 36830 11040 36864
rect 10984 36796 11040 36830
rect 10984 36762 10995 36796
rect 11029 36762 11040 36796
rect 10984 36728 11040 36762
rect 10984 36694 10995 36728
rect 11029 36694 11040 36728
rect 10984 36660 11040 36694
rect 10984 36626 10995 36660
rect 11029 36626 11040 36660
rect 10984 36592 11040 36626
rect 10984 36558 10995 36592
rect 11029 36558 11040 36592
rect 10984 36524 11040 36558
rect 10984 36490 10995 36524
rect 11029 36490 11040 36524
rect 10984 36456 11040 36490
rect 10984 36422 10995 36456
rect 11029 36422 11040 36456
rect 10984 36388 11040 36422
rect 10984 36354 10995 36388
rect 11029 36354 11040 36388
rect 10984 36320 11040 36354
rect 10984 36286 10995 36320
rect 11029 36286 11040 36320
rect 10984 36252 11040 36286
rect 10984 36218 10995 36252
rect 11029 36218 11040 36252
rect 10984 36184 11040 36218
rect 10984 36150 10995 36184
rect 11029 36150 11040 36184
rect 10984 36116 11040 36150
rect 10984 36082 10995 36116
rect 11029 36082 11040 36116
rect 10984 36036 11040 36082
rect 11640 37340 11696 37386
rect 11640 37306 11651 37340
rect 11685 37306 11696 37340
rect 11640 37272 11696 37306
rect 11640 37238 11651 37272
rect 11685 37238 11696 37272
rect 11640 37204 11696 37238
rect 11640 37170 11651 37204
rect 11685 37170 11696 37204
rect 11640 37136 11696 37170
rect 11640 37102 11651 37136
rect 11685 37102 11696 37136
rect 11640 37068 11696 37102
rect 11640 37034 11651 37068
rect 11685 37034 11696 37068
rect 11640 37000 11696 37034
rect 11640 36966 11651 37000
rect 11685 36966 11696 37000
rect 11640 36932 11696 36966
rect 11640 36898 11651 36932
rect 11685 36898 11696 36932
rect 11640 36864 11696 36898
rect 11640 36830 11651 36864
rect 11685 36830 11696 36864
rect 11640 36796 11696 36830
rect 11640 36762 11651 36796
rect 11685 36762 11696 36796
rect 11640 36728 11696 36762
rect 11640 36694 11651 36728
rect 11685 36694 11696 36728
rect 11640 36660 11696 36694
rect 11640 36626 11651 36660
rect 11685 36626 11696 36660
rect 11640 36592 11696 36626
rect 11640 36558 11651 36592
rect 11685 36558 11696 36592
rect 11640 36524 11696 36558
rect 11640 36490 11651 36524
rect 11685 36490 11696 36524
rect 11640 36456 11696 36490
rect 11640 36422 11651 36456
rect 11685 36422 11696 36456
rect 11640 36388 11696 36422
rect 11640 36354 11651 36388
rect 11685 36354 11696 36388
rect 11640 36320 11696 36354
rect 11640 36286 11651 36320
rect 11685 36286 11696 36320
rect 11640 36252 11696 36286
rect 11640 36218 11651 36252
rect 11685 36218 11696 36252
rect 11640 36184 11696 36218
rect 11640 36150 11651 36184
rect 11685 36150 11696 36184
rect 11640 36116 11696 36150
rect 11640 36082 11651 36116
rect 11685 36082 11696 36116
rect 11640 36036 11696 36082
rect 12296 37340 12352 37386
rect 12296 37306 12307 37340
rect 12341 37306 12352 37340
rect 12296 37272 12352 37306
rect 12296 37238 12307 37272
rect 12341 37238 12352 37272
rect 12296 37204 12352 37238
rect 12296 37170 12307 37204
rect 12341 37170 12352 37204
rect 12296 37136 12352 37170
rect 12296 37102 12307 37136
rect 12341 37102 12352 37136
rect 12296 37068 12352 37102
rect 12296 37034 12307 37068
rect 12341 37034 12352 37068
rect 12296 37000 12352 37034
rect 12296 36966 12307 37000
rect 12341 36966 12352 37000
rect 12296 36932 12352 36966
rect 12296 36898 12307 36932
rect 12341 36898 12352 36932
rect 12296 36864 12352 36898
rect 12296 36830 12307 36864
rect 12341 36830 12352 36864
rect 12296 36796 12352 36830
rect 12296 36762 12307 36796
rect 12341 36762 12352 36796
rect 12296 36728 12352 36762
rect 12296 36694 12307 36728
rect 12341 36694 12352 36728
rect 12296 36660 12352 36694
rect 12296 36626 12307 36660
rect 12341 36626 12352 36660
rect 12296 36592 12352 36626
rect 12296 36558 12307 36592
rect 12341 36558 12352 36592
rect 12296 36524 12352 36558
rect 12296 36490 12307 36524
rect 12341 36490 12352 36524
rect 12296 36456 12352 36490
rect 12296 36422 12307 36456
rect 12341 36422 12352 36456
rect 12296 36388 12352 36422
rect 12296 36354 12307 36388
rect 12341 36354 12352 36388
rect 12296 36320 12352 36354
rect 12296 36286 12307 36320
rect 12341 36286 12352 36320
rect 12296 36252 12352 36286
rect 12296 36218 12307 36252
rect 12341 36218 12352 36252
rect 12296 36184 12352 36218
rect 12296 36150 12307 36184
rect 12341 36150 12352 36184
rect 12296 36116 12352 36150
rect 12296 36082 12307 36116
rect 12341 36082 12352 36116
rect 12296 36036 12352 36082
rect 12952 37340 13008 37386
rect 12952 37306 12963 37340
rect 12997 37306 13008 37340
rect 12952 37272 13008 37306
rect 12952 37238 12963 37272
rect 12997 37238 13008 37272
rect 12952 37204 13008 37238
rect 12952 37170 12963 37204
rect 12997 37170 13008 37204
rect 12952 37136 13008 37170
rect 12952 37102 12963 37136
rect 12997 37102 13008 37136
rect 12952 37068 13008 37102
rect 12952 37034 12963 37068
rect 12997 37034 13008 37068
rect 12952 37000 13008 37034
rect 12952 36966 12963 37000
rect 12997 36966 13008 37000
rect 12952 36932 13008 36966
rect 12952 36898 12963 36932
rect 12997 36898 13008 36932
rect 12952 36864 13008 36898
rect 12952 36830 12963 36864
rect 12997 36830 13008 36864
rect 12952 36796 13008 36830
rect 12952 36762 12963 36796
rect 12997 36762 13008 36796
rect 12952 36728 13008 36762
rect 12952 36694 12963 36728
rect 12997 36694 13008 36728
rect 12952 36660 13008 36694
rect 12952 36626 12963 36660
rect 12997 36626 13008 36660
rect 12952 36592 13008 36626
rect 12952 36558 12963 36592
rect 12997 36558 13008 36592
rect 12952 36524 13008 36558
rect 12952 36490 12963 36524
rect 12997 36490 13008 36524
rect 12952 36456 13008 36490
rect 12952 36422 12963 36456
rect 12997 36422 13008 36456
rect 12952 36388 13008 36422
rect 12952 36354 12963 36388
rect 12997 36354 13008 36388
rect 12952 36320 13008 36354
rect 12952 36286 12963 36320
rect 12997 36286 13008 36320
rect 12952 36252 13008 36286
rect 12952 36218 12963 36252
rect 12997 36218 13008 36252
rect 12952 36184 13008 36218
rect 12952 36150 12963 36184
rect 12997 36150 13008 36184
rect 12952 36116 13008 36150
rect 12952 36082 12963 36116
rect 12997 36082 13008 36116
rect 12952 36036 13008 36082
rect 13608 37340 13664 37386
rect 13608 37306 13619 37340
rect 13653 37306 13664 37340
rect 13608 37272 13664 37306
rect 13608 37238 13619 37272
rect 13653 37238 13664 37272
rect 13608 37204 13664 37238
rect 13608 37170 13619 37204
rect 13653 37170 13664 37204
rect 13608 37136 13664 37170
rect 13608 37102 13619 37136
rect 13653 37102 13664 37136
rect 13608 37068 13664 37102
rect 13608 37034 13619 37068
rect 13653 37034 13664 37068
rect 13608 37000 13664 37034
rect 13608 36966 13619 37000
rect 13653 36966 13664 37000
rect 13608 36932 13664 36966
rect 13608 36898 13619 36932
rect 13653 36898 13664 36932
rect 13608 36864 13664 36898
rect 13608 36830 13619 36864
rect 13653 36830 13664 36864
rect 13608 36796 13664 36830
rect 13608 36762 13619 36796
rect 13653 36762 13664 36796
rect 13608 36728 13664 36762
rect 13608 36694 13619 36728
rect 13653 36694 13664 36728
rect 13608 36660 13664 36694
rect 13608 36626 13619 36660
rect 13653 36626 13664 36660
rect 13608 36592 13664 36626
rect 13608 36558 13619 36592
rect 13653 36558 13664 36592
rect 13608 36524 13664 36558
rect 13608 36490 13619 36524
rect 13653 36490 13664 36524
rect 13608 36456 13664 36490
rect 13608 36422 13619 36456
rect 13653 36422 13664 36456
rect 13608 36388 13664 36422
rect 13608 36354 13619 36388
rect 13653 36354 13664 36388
rect 13608 36320 13664 36354
rect 13608 36286 13619 36320
rect 13653 36286 13664 36320
rect 13608 36252 13664 36286
rect 13608 36218 13619 36252
rect 13653 36218 13664 36252
rect 13608 36184 13664 36218
rect 13608 36150 13619 36184
rect 13653 36150 13664 36184
rect 13608 36116 13664 36150
rect 13608 36082 13619 36116
rect 13653 36082 13664 36116
rect 13608 36036 13664 36082
rect 14264 37340 14317 37386
rect 14264 37306 14275 37340
rect 14309 37306 14317 37340
rect 14264 37272 14317 37306
rect 14264 37238 14275 37272
rect 14309 37238 14317 37272
rect 14264 37204 14317 37238
rect 14264 37170 14275 37204
rect 14309 37170 14317 37204
rect 14264 37136 14317 37170
rect 14264 37102 14275 37136
rect 14309 37102 14317 37136
rect 14264 37068 14317 37102
rect 14264 37034 14275 37068
rect 14309 37034 14317 37068
rect 14264 37000 14317 37034
rect 14264 36966 14275 37000
rect 14309 36966 14317 37000
rect 14264 36932 14317 36966
rect 14264 36898 14275 36932
rect 14309 36898 14317 36932
rect 14264 36864 14317 36898
rect 14264 36830 14275 36864
rect 14309 36830 14317 36864
rect 14264 36796 14317 36830
rect 14264 36762 14275 36796
rect 14309 36762 14317 36796
rect 14264 36728 14317 36762
rect 14264 36694 14275 36728
rect 14309 36694 14317 36728
rect 14264 36660 14317 36694
rect 14264 36626 14275 36660
rect 14309 36626 14317 36660
rect 14264 36592 14317 36626
rect 14264 36558 14275 36592
rect 14309 36558 14317 36592
rect 14264 36524 14317 36558
rect 14264 36490 14275 36524
rect 14309 36490 14317 36524
rect 14264 36456 14317 36490
rect 14264 36422 14275 36456
rect 14309 36422 14317 36456
rect 14264 36388 14317 36422
rect 14264 36354 14275 36388
rect 14309 36354 14317 36388
rect 14264 36320 14317 36354
rect 14264 36286 14275 36320
rect 14309 36286 14317 36320
rect 14264 36252 14317 36286
rect 14264 36218 14275 36252
rect 14309 36218 14317 36252
rect 14264 36184 14317 36218
rect 14264 36150 14275 36184
rect 14309 36150 14317 36184
rect 14264 36116 14317 36150
rect 14264 36082 14275 36116
rect 14309 36082 14317 36116
rect 14264 36036 14317 36082
rect 9569 35918 9622 35964
rect 9569 35884 9577 35918
rect 9611 35884 9622 35918
rect 9569 35850 9622 35884
rect 9569 35816 9577 35850
rect 9611 35816 9622 35850
rect 9569 35782 9622 35816
rect 9569 35748 9577 35782
rect 9611 35748 9622 35782
rect 9569 35714 9622 35748
rect 9569 35680 9577 35714
rect 9611 35680 9622 35714
rect 9569 35646 9622 35680
rect 9569 35612 9577 35646
rect 9611 35612 9622 35646
rect 9569 35578 9622 35612
rect 9569 35544 9577 35578
rect 9611 35544 9622 35578
rect 9569 35510 9622 35544
rect 9569 35476 9577 35510
rect 9611 35476 9622 35510
rect 9569 35442 9622 35476
rect 9569 35408 9577 35442
rect 9611 35408 9622 35442
rect 9569 35374 9622 35408
rect 9569 35340 9577 35374
rect 9611 35340 9622 35374
rect 9569 35306 9622 35340
rect 9569 35272 9577 35306
rect 9611 35272 9622 35306
rect 9569 35238 9622 35272
rect 9569 35204 9577 35238
rect 9611 35204 9622 35238
rect 9569 35170 9622 35204
rect 9569 35136 9577 35170
rect 9611 35136 9622 35170
rect 9569 35102 9622 35136
rect 9569 35068 9577 35102
rect 9611 35068 9622 35102
rect 9569 35034 9622 35068
rect 9569 35000 9577 35034
rect 9611 35000 9622 35034
rect 9569 34966 9622 35000
rect 9569 34932 9577 34966
rect 9611 34932 9622 34966
rect 9569 34898 9622 34932
rect 9569 34864 9577 34898
rect 9611 34864 9622 34898
rect 9569 34830 9622 34864
rect 9569 34796 9577 34830
rect 9611 34796 9622 34830
rect 9569 34762 9622 34796
rect 9569 34728 9577 34762
rect 9611 34728 9622 34762
rect 9569 34694 9622 34728
rect 9569 34660 9577 34694
rect 9611 34660 9622 34694
rect 9569 34614 9622 34660
rect 10222 35918 10275 35964
rect 10222 35884 10233 35918
rect 10267 35884 10275 35918
rect 10222 35850 10275 35884
rect 10222 35816 10233 35850
rect 10267 35816 10275 35850
rect 10222 35782 10275 35816
rect 10222 35748 10233 35782
rect 10267 35748 10275 35782
rect 10222 35714 10275 35748
rect 10222 35680 10233 35714
rect 10267 35680 10275 35714
rect 10222 35646 10275 35680
rect 10222 35612 10233 35646
rect 10267 35612 10275 35646
rect 10222 35578 10275 35612
rect 10222 35544 10233 35578
rect 10267 35544 10275 35578
rect 10222 35510 10275 35544
rect 10222 35476 10233 35510
rect 10267 35476 10275 35510
rect 10222 35442 10275 35476
rect 10222 35408 10233 35442
rect 10267 35408 10275 35442
rect 10222 35374 10275 35408
rect 10222 35340 10233 35374
rect 10267 35340 10275 35374
rect 10222 35306 10275 35340
rect 10222 35272 10233 35306
rect 10267 35272 10275 35306
rect 10222 35238 10275 35272
rect 10222 35204 10233 35238
rect 10267 35204 10275 35238
rect 10222 35170 10275 35204
rect 10222 35136 10233 35170
rect 10267 35136 10275 35170
rect 10222 35102 10275 35136
rect 10222 35068 10233 35102
rect 10267 35068 10275 35102
rect 10222 35034 10275 35068
rect 10222 35000 10233 35034
rect 10267 35000 10275 35034
rect 10222 34966 10275 35000
rect 10222 34932 10233 34966
rect 10267 34932 10275 34966
rect 10222 34898 10275 34932
rect 10222 34864 10233 34898
rect 10267 34864 10275 34898
rect 10222 34830 10275 34864
rect 10222 34796 10233 34830
rect 10267 34796 10275 34830
rect 10222 34762 10275 34796
rect 10222 34728 10233 34762
rect 10267 34728 10275 34762
rect 10222 34694 10275 34728
rect 10222 34660 10233 34694
rect 10267 34660 10275 34694
rect 10222 34614 10275 34660
rect 10331 35918 10384 35964
rect 10331 35884 10339 35918
rect 10373 35884 10384 35918
rect 10331 35850 10384 35884
rect 10331 35816 10339 35850
rect 10373 35816 10384 35850
rect 10331 35782 10384 35816
rect 10331 35748 10339 35782
rect 10373 35748 10384 35782
rect 10331 35714 10384 35748
rect 10331 35680 10339 35714
rect 10373 35680 10384 35714
rect 10331 35646 10384 35680
rect 10331 35612 10339 35646
rect 10373 35612 10384 35646
rect 10331 35578 10384 35612
rect 10331 35544 10339 35578
rect 10373 35544 10384 35578
rect 10331 35510 10384 35544
rect 10331 35476 10339 35510
rect 10373 35476 10384 35510
rect 10331 35442 10384 35476
rect 10331 35408 10339 35442
rect 10373 35408 10384 35442
rect 10331 35374 10384 35408
rect 10331 35340 10339 35374
rect 10373 35340 10384 35374
rect 10331 35306 10384 35340
rect 10331 35272 10339 35306
rect 10373 35272 10384 35306
rect 10331 35238 10384 35272
rect 10331 35204 10339 35238
rect 10373 35204 10384 35238
rect 10331 35170 10384 35204
rect 10331 35136 10339 35170
rect 10373 35136 10384 35170
rect 10331 35102 10384 35136
rect 10331 35068 10339 35102
rect 10373 35068 10384 35102
rect 10331 35034 10384 35068
rect 10331 35000 10339 35034
rect 10373 35000 10384 35034
rect 10331 34966 10384 35000
rect 10331 34932 10339 34966
rect 10373 34932 10384 34966
rect 10331 34898 10384 34932
rect 10331 34864 10339 34898
rect 10373 34864 10384 34898
rect 10331 34830 10384 34864
rect 10331 34796 10339 34830
rect 10373 34796 10384 34830
rect 10331 34762 10384 34796
rect 10331 34728 10339 34762
rect 10373 34728 10384 34762
rect 10331 34694 10384 34728
rect 10331 34660 10339 34694
rect 10373 34660 10384 34694
rect 10331 34614 10384 34660
rect 10984 35918 11040 35964
rect 10984 35884 10995 35918
rect 11029 35884 11040 35918
rect 10984 35850 11040 35884
rect 10984 35816 10995 35850
rect 11029 35816 11040 35850
rect 10984 35782 11040 35816
rect 10984 35748 10995 35782
rect 11029 35748 11040 35782
rect 10984 35714 11040 35748
rect 10984 35680 10995 35714
rect 11029 35680 11040 35714
rect 10984 35646 11040 35680
rect 10984 35612 10995 35646
rect 11029 35612 11040 35646
rect 10984 35578 11040 35612
rect 10984 35544 10995 35578
rect 11029 35544 11040 35578
rect 10984 35510 11040 35544
rect 10984 35476 10995 35510
rect 11029 35476 11040 35510
rect 10984 35442 11040 35476
rect 10984 35408 10995 35442
rect 11029 35408 11040 35442
rect 10984 35374 11040 35408
rect 10984 35340 10995 35374
rect 11029 35340 11040 35374
rect 10984 35306 11040 35340
rect 10984 35272 10995 35306
rect 11029 35272 11040 35306
rect 10984 35238 11040 35272
rect 10984 35204 10995 35238
rect 11029 35204 11040 35238
rect 10984 35170 11040 35204
rect 10984 35136 10995 35170
rect 11029 35136 11040 35170
rect 10984 35102 11040 35136
rect 10984 35068 10995 35102
rect 11029 35068 11040 35102
rect 10984 35034 11040 35068
rect 10984 35000 10995 35034
rect 11029 35000 11040 35034
rect 10984 34966 11040 35000
rect 10984 34932 10995 34966
rect 11029 34932 11040 34966
rect 10984 34898 11040 34932
rect 10984 34864 10995 34898
rect 11029 34864 11040 34898
rect 10984 34830 11040 34864
rect 10984 34796 10995 34830
rect 11029 34796 11040 34830
rect 10984 34762 11040 34796
rect 10984 34728 10995 34762
rect 11029 34728 11040 34762
rect 10984 34694 11040 34728
rect 10984 34660 10995 34694
rect 11029 34660 11040 34694
rect 10984 34614 11040 34660
rect 11640 35918 11696 35964
rect 11640 35884 11651 35918
rect 11685 35884 11696 35918
rect 11640 35850 11696 35884
rect 11640 35816 11651 35850
rect 11685 35816 11696 35850
rect 11640 35782 11696 35816
rect 11640 35748 11651 35782
rect 11685 35748 11696 35782
rect 11640 35714 11696 35748
rect 11640 35680 11651 35714
rect 11685 35680 11696 35714
rect 11640 35646 11696 35680
rect 11640 35612 11651 35646
rect 11685 35612 11696 35646
rect 11640 35578 11696 35612
rect 11640 35544 11651 35578
rect 11685 35544 11696 35578
rect 11640 35510 11696 35544
rect 11640 35476 11651 35510
rect 11685 35476 11696 35510
rect 11640 35442 11696 35476
rect 11640 35408 11651 35442
rect 11685 35408 11696 35442
rect 11640 35374 11696 35408
rect 11640 35340 11651 35374
rect 11685 35340 11696 35374
rect 11640 35306 11696 35340
rect 11640 35272 11651 35306
rect 11685 35272 11696 35306
rect 11640 35238 11696 35272
rect 11640 35204 11651 35238
rect 11685 35204 11696 35238
rect 11640 35170 11696 35204
rect 11640 35136 11651 35170
rect 11685 35136 11696 35170
rect 11640 35102 11696 35136
rect 11640 35068 11651 35102
rect 11685 35068 11696 35102
rect 11640 35034 11696 35068
rect 11640 35000 11651 35034
rect 11685 35000 11696 35034
rect 11640 34966 11696 35000
rect 11640 34932 11651 34966
rect 11685 34932 11696 34966
rect 11640 34898 11696 34932
rect 11640 34864 11651 34898
rect 11685 34864 11696 34898
rect 11640 34830 11696 34864
rect 11640 34796 11651 34830
rect 11685 34796 11696 34830
rect 11640 34762 11696 34796
rect 11640 34728 11651 34762
rect 11685 34728 11696 34762
rect 11640 34694 11696 34728
rect 11640 34660 11651 34694
rect 11685 34660 11696 34694
rect 11640 34614 11696 34660
rect 12296 35918 12352 35964
rect 12296 35884 12307 35918
rect 12341 35884 12352 35918
rect 12296 35850 12352 35884
rect 12296 35816 12307 35850
rect 12341 35816 12352 35850
rect 12296 35782 12352 35816
rect 12296 35748 12307 35782
rect 12341 35748 12352 35782
rect 12296 35714 12352 35748
rect 12296 35680 12307 35714
rect 12341 35680 12352 35714
rect 12296 35646 12352 35680
rect 12296 35612 12307 35646
rect 12341 35612 12352 35646
rect 12296 35578 12352 35612
rect 12296 35544 12307 35578
rect 12341 35544 12352 35578
rect 12296 35510 12352 35544
rect 12296 35476 12307 35510
rect 12341 35476 12352 35510
rect 12296 35442 12352 35476
rect 12296 35408 12307 35442
rect 12341 35408 12352 35442
rect 12296 35374 12352 35408
rect 12296 35340 12307 35374
rect 12341 35340 12352 35374
rect 12296 35306 12352 35340
rect 12296 35272 12307 35306
rect 12341 35272 12352 35306
rect 12296 35238 12352 35272
rect 12296 35204 12307 35238
rect 12341 35204 12352 35238
rect 12296 35170 12352 35204
rect 12296 35136 12307 35170
rect 12341 35136 12352 35170
rect 12296 35102 12352 35136
rect 12296 35068 12307 35102
rect 12341 35068 12352 35102
rect 12296 35034 12352 35068
rect 12296 35000 12307 35034
rect 12341 35000 12352 35034
rect 12296 34966 12352 35000
rect 12296 34932 12307 34966
rect 12341 34932 12352 34966
rect 12296 34898 12352 34932
rect 12296 34864 12307 34898
rect 12341 34864 12352 34898
rect 12296 34830 12352 34864
rect 12296 34796 12307 34830
rect 12341 34796 12352 34830
rect 12296 34762 12352 34796
rect 12296 34728 12307 34762
rect 12341 34728 12352 34762
rect 12296 34694 12352 34728
rect 12296 34660 12307 34694
rect 12341 34660 12352 34694
rect 12296 34614 12352 34660
rect 12952 35918 13008 35964
rect 12952 35884 12963 35918
rect 12997 35884 13008 35918
rect 12952 35850 13008 35884
rect 12952 35816 12963 35850
rect 12997 35816 13008 35850
rect 12952 35782 13008 35816
rect 12952 35748 12963 35782
rect 12997 35748 13008 35782
rect 12952 35714 13008 35748
rect 12952 35680 12963 35714
rect 12997 35680 13008 35714
rect 12952 35646 13008 35680
rect 12952 35612 12963 35646
rect 12997 35612 13008 35646
rect 12952 35578 13008 35612
rect 12952 35544 12963 35578
rect 12997 35544 13008 35578
rect 12952 35510 13008 35544
rect 12952 35476 12963 35510
rect 12997 35476 13008 35510
rect 12952 35442 13008 35476
rect 12952 35408 12963 35442
rect 12997 35408 13008 35442
rect 12952 35374 13008 35408
rect 12952 35340 12963 35374
rect 12997 35340 13008 35374
rect 12952 35306 13008 35340
rect 12952 35272 12963 35306
rect 12997 35272 13008 35306
rect 12952 35238 13008 35272
rect 12952 35204 12963 35238
rect 12997 35204 13008 35238
rect 12952 35170 13008 35204
rect 12952 35136 12963 35170
rect 12997 35136 13008 35170
rect 12952 35102 13008 35136
rect 12952 35068 12963 35102
rect 12997 35068 13008 35102
rect 12952 35034 13008 35068
rect 12952 35000 12963 35034
rect 12997 35000 13008 35034
rect 12952 34966 13008 35000
rect 12952 34932 12963 34966
rect 12997 34932 13008 34966
rect 12952 34898 13008 34932
rect 12952 34864 12963 34898
rect 12997 34864 13008 34898
rect 12952 34830 13008 34864
rect 12952 34796 12963 34830
rect 12997 34796 13008 34830
rect 12952 34762 13008 34796
rect 12952 34728 12963 34762
rect 12997 34728 13008 34762
rect 12952 34694 13008 34728
rect 12952 34660 12963 34694
rect 12997 34660 13008 34694
rect 12952 34614 13008 34660
rect 13608 35918 13664 35964
rect 13608 35884 13619 35918
rect 13653 35884 13664 35918
rect 13608 35850 13664 35884
rect 13608 35816 13619 35850
rect 13653 35816 13664 35850
rect 13608 35782 13664 35816
rect 13608 35748 13619 35782
rect 13653 35748 13664 35782
rect 13608 35714 13664 35748
rect 13608 35680 13619 35714
rect 13653 35680 13664 35714
rect 13608 35646 13664 35680
rect 13608 35612 13619 35646
rect 13653 35612 13664 35646
rect 13608 35578 13664 35612
rect 13608 35544 13619 35578
rect 13653 35544 13664 35578
rect 13608 35510 13664 35544
rect 13608 35476 13619 35510
rect 13653 35476 13664 35510
rect 13608 35442 13664 35476
rect 13608 35408 13619 35442
rect 13653 35408 13664 35442
rect 13608 35374 13664 35408
rect 13608 35340 13619 35374
rect 13653 35340 13664 35374
rect 13608 35306 13664 35340
rect 13608 35272 13619 35306
rect 13653 35272 13664 35306
rect 13608 35238 13664 35272
rect 13608 35204 13619 35238
rect 13653 35204 13664 35238
rect 13608 35170 13664 35204
rect 13608 35136 13619 35170
rect 13653 35136 13664 35170
rect 13608 35102 13664 35136
rect 13608 35068 13619 35102
rect 13653 35068 13664 35102
rect 13608 35034 13664 35068
rect 13608 35000 13619 35034
rect 13653 35000 13664 35034
rect 13608 34966 13664 35000
rect 13608 34932 13619 34966
rect 13653 34932 13664 34966
rect 13608 34898 13664 34932
rect 13608 34864 13619 34898
rect 13653 34864 13664 34898
rect 13608 34830 13664 34864
rect 13608 34796 13619 34830
rect 13653 34796 13664 34830
rect 13608 34762 13664 34796
rect 13608 34728 13619 34762
rect 13653 34728 13664 34762
rect 13608 34694 13664 34728
rect 13608 34660 13619 34694
rect 13653 34660 13664 34694
rect 13608 34614 13664 34660
rect 14264 35918 14317 35964
rect 14264 35884 14275 35918
rect 14309 35884 14317 35918
rect 14264 35850 14317 35884
rect 14264 35816 14275 35850
rect 14309 35816 14317 35850
rect 14264 35782 14317 35816
rect 14264 35748 14275 35782
rect 14309 35748 14317 35782
rect 14264 35714 14317 35748
rect 14264 35680 14275 35714
rect 14309 35680 14317 35714
rect 14264 35646 14317 35680
rect 14264 35612 14275 35646
rect 14309 35612 14317 35646
rect 14264 35578 14317 35612
rect 14264 35544 14275 35578
rect 14309 35544 14317 35578
rect 14264 35510 14317 35544
rect 14264 35476 14275 35510
rect 14309 35476 14317 35510
rect 14264 35442 14317 35476
rect 14264 35408 14275 35442
rect 14309 35408 14317 35442
rect 14264 35374 14317 35408
rect 14264 35340 14275 35374
rect 14309 35340 14317 35374
rect 14264 35306 14317 35340
rect 14264 35272 14275 35306
rect 14309 35272 14317 35306
rect 14264 35238 14317 35272
rect 14264 35204 14275 35238
rect 14309 35204 14317 35238
rect 14264 35170 14317 35204
rect 14264 35136 14275 35170
rect 14309 35136 14317 35170
rect 14264 35102 14317 35136
rect 14264 35068 14275 35102
rect 14309 35068 14317 35102
rect 14264 35034 14317 35068
rect 14264 35000 14275 35034
rect 14309 35000 14317 35034
rect 14264 34966 14317 35000
rect 14264 34932 14275 34966
rect 14309 34932 14317 34966
rect 14264 34898 14317 34932
rect 14264 34864 14275 34898
rect 14309 34864 14317 34898
rect 14264 34830 14317 34864
rect 14264 34796 14275 34830
rect 14309 34796 14317 34830
rect 14264 34762 14317 34796
rect 14264 34728 14275 34762
rect 14309 34728 14317 34762
rect 14264 34694 14317 34728
rect 14264 34660 14275 34694
rect 14309 34660 14317 34694
rect 14264 34614 14317 34660
rect 19087 37322 19132 37368
rect 19121 37288 19132 37322
rect 19087 37254 19132 37288
rect 19121 37220 19132 37254
rect 19087 37186 19132 37220
rect 19121 37152 19132 37186
rect 19087 37118 19132 37152
rect 19121 37084 19132 37118
rect 19087 37050 19132 37084
rect 19121 37016 19132 37050
rect 19087 36982 19132 37016
rect 19121 36948 19132 36982
rect 19087 36914 19132 36948
rect 19121 36880 19132 36914
rect 19087 36846 19132 36880
rect 19121 36812 19132 36846
rect 19087 36778 19132 36812
rect 19121 36744 19132 36778
rect 19087 36710 19132 36744
rect 19121 36676 19132 36710
rect 19087 36642 19132 36676
rect 19121 36608 19132 36642
rect 19087 36574 19132 36608
rect 19121 36540 19132 36574
rect 19087 36506 19132 36540
rect 19121 36472 19132 36506
rect 19087 36438 19132 36472
rect 19121 36404 19132 36438
rect 19087 36370 19132 36404
rect 19121 36336 19132 36370
rect 19087 36302 19132 36336
rect 19121 36268 19132 36302
rect 19087 36234 19132 36268
rect 19121 36200 19132 36234
rect 19087 36166 19132 36200
rect 19121 36132 19132 36166
rect 19087 36098 19132 36132
rect 19121 36064 19132 36098
rect 19087 36018 19132 36064
rect 19732 37322 19788 37368
rect 19732 37288 19743 37322
rect 19777 37288 19788 37322
rect 19732 37254 19788 37288
rect 19732 37220 19743 37254
rect 19777 37220 19788 37254
rect 19732 37186 19788 37220
rect 19732 37152 19743 37186
rect 19777 37152 19788 37186
rect 19732 37118 19788 37152
rect 19732 37084 19743 37118
rect 19777 37084 19788 37118
rect 19732 37050 19788 37084
rect 19732 37016 19743 37050
rect 19777 37016 19788 37050
rect 19732 36982 19788 37016
rect 19732 36948 19743 36982
rect 19777 36948 19788 36982
rect 19732 36914 19788 36948
rect 19732 36880 19743 36914
rect 19777 36880 19788 36914
rect 19732 36846 19788 36880
rect 19732 36812 19743 36846
rect 19777 36812 19788 36846
rect 19732 36778 19788 36812
rect 19732 36744 19743 36778
rect 19777 36744 19788 36778
rect 19732 36710 19788 36744
rect 19732 36676 19743 36710
rect 19777 36676 19788 36710
rect 19732 36642 19788 36676
rect 19732 36608 19743 36642
rect 19777 36608 19788 36642
rect 19732 36574 19788 36608
rect 19732 36540 19743 36574
rect 19777 36540 19788 36574
rect 19732 36506 19788 36540
rect 19732 36472 19743 36506
rect 19777 36472 19788 36506
rect 19732 36438 19788 36472
rect 19732 36404 19743 36438
rect 19777 36404 19788 36438
rect 19732 36370 19788 36404
rect 19732 36336 19743 36370
rect 19777 36336 19788 36370
rect 19732 36302 19788 36336
rect 19732 36268 19743 36302
rect 19777 36268 19788 36302
rect 19732 36234 19788 36268
rect 19732 36200 19743 36234
rect 19777 36200 19788 36234
rect 19732 36166 19788 36200
rect 19732 36132 19743 36166
rect 19777 36132 19788 36166
rect 19732 36098 19788 36132
rect 19732 36064 19743 36098
rect 19777 36064 19788 36098
rect 19732 36018 19788 36064
rect 20388 37322 20444 37368
rect 20388 37288 20399 37322
rect 20433 37288 20444 37322
rect 20388 37254 20444 37288
rect 20388 37220 20399 37254
rect 20433 37220 20444 37254
rect 20388 37186 20444 37220
rect 20388 37152 20399 37186
rect 20433 37152 20444 37186
rect 20388 37118 20444 37152
rect 20388 37084 20399 37118
rect 20433 37084 20444 37118
rect 20388 37050 20444 37084
rect 20388 37016 20399 37050
rect 20433 37016 20444 37050
rect 20388 36982 20444 37016
rect 20388 36948 20399 36982
rect 20433 36948 20444 36982
rect 20388 36914 20444 36948
rect 20388 36880 20399 36914
rect 20433 36880 20444 36914
rect 20388 36846 20444 36880
rect 20388 36812 20399 36846
rect 20433 36812 20444 36846
rect 20388 36778 20444 36812
rect 20388 36744 20399 36778
rect 20433 36744 20444 36778
rect 20388 36710 20444 36744
rect 20388 36676 20399 36710
rect 20433 36676 20444 36710
rect 20388 36642 20444 36676
rect 20388 36608 20399 36642
rect 20433 36608 20444 36642
rect 20388 36574 20444 36608
rect 20388 36540 20399 36574
rect 20433 36540 20444 36574
rect 20388 36506 20444 36540
rect 20388 36472 20399 36506
rect 20433 36472 20444 36506
rect 20388 36438 20444 36472
rect 20388 36404 20399 36438
rect 20433 36404 20444 36438
rect 20388 36370 20444 36404
rect 20388 36336 20399 36370
rect 20433 36336 20444 36370
rect 20388 36302 20444 36336
rect 20388 36268 20399 36302
rect 20433 36268 20444 36302
rect 20388 36234 20444 36268
rect 20388 36200 20399 36234
rect 20433 36200 20444 36234
rect 20388 36166 20444 36200
rect 20388 36132 20399 36166
rect 20433 36132 20444 36166
rect 20388 36098 20444 36132
rect 20388 36064 20399 36098
rect 20433 36064 20444 36098
rect 20388 36018 20444 36064
rect 21044 37322 21100 37368
rect 21044 37288 21055 37322
rect 21089 37288 21100 37322
rect 21044 37254 21100 37288
rect 21044 37220 21055 37254
rect 21089 37220 21100 37254
rect 21044 37186 21100 37220
rect 21044 37152 21055 37186
rect 21089 37152 21100 37186
rect 21044 37118 21100 37152
rect 21044 37084 21055 37118
rect 21089 37084 21100 37118
rect 21044 37050 21100 37084
rect 21044 37016 21055 37050
rect 21089 37016 21100 37050
rect 21044 36982 21100 37016
rect 21044 36948 21055 36982
rect 21089 36948 21100 36982
rect 21044 36914 21100 36948
rect 21044 36880 21055 36914
rect 21089 36880 21100 36914
rect 21044 36846 21100 36880
rect 21044 36812 21055 36846
rect 21089 36812 21100 36846
rect 21044 36778 21100 36812
rect 21044 36744 21055 36778
rect 21089 36744 21100 36778
rect 21044 36710 21100 36744
rect 21044 36676 21055 36710
rect 21089 36676 21100 36710
rect 21044 36642 21100 36676
rect 21044 36608 21055 36642
rect 21089 36608 21100 36642
rect 21044 36574 21100 36608
rect 21044 36540 21055 36574
rect 21089 36540 21100 36574
rect 21044 36506 21100 36540
rect 21044 36472 21055 36506
rect 21089 36472 21100 36506
rect 21044 36438 21100 36472
rect 21044 36404 21055 36438
rect 21089 36404 21100 36438
rect 21044 36370 21100 36404
rect 21044 36336 21055 36370
rect 21089 36336 21100 36370
rect 21044 36302 21100 36336
rect 21044 36268 21055 36302
rect 21089 36268 21100 36302
rect 21044 36234 21100 36268
rect 21044 36200 21055 36234
rect 21089 36200 21100 36234
rect 21044 36166 21100 36200
rect 21044 36132 21055 36166
rect 21089 36132 21100 36166
rect 21044 36098 21100 36132
rect 21044 36064 21055 36098
rect 21089 36064 21100 36098
rect 21044 36018 21100 36064
rect 21700 37322 21756 37368
rect 21700 37288 21711 37322
rect 21745 37288 21756 37322
rect 21700 37254 21756 37288
rect 21700 37220 21711 37254
rect 21745 37220 21756 37254
rect 21700 37186 21756 37220
rect 21700 37152 21711 37186
rect 21745 37152 21756 37186
rect 21700 37118 21756 37152
rect 21700 37084 21711 37118
rect 21745 37084 21756 37118
rect 21700 37050 21756 37084
rect 21700 37016 21711 37050
rect 21745 37016 21756 37050
rect 21700 36982 21756 37016
rect 21700 36948 21711 36982
rect 21745 36948 21756 36982
rect 21700 36914 21756 36948
rect 21700 36880 21711 36914
rect 21745 36880 21756 36914
rect 21700 36846 21756 36880
rect 21700 36812 21711 36846
rect 21745 36812 21756 36846
rect 21700 36778 21756 36812
rect 21700 36744 21711 36778
rect 21745 36744 21756 36778
rect 21700 36710 21756 36744
rect 21700 36676 21711 36710
rect 21745 36676 21756 36710
rect 21700 36642 21756 36676
rect 21700 36608 21711 36642
rect 21745 36608 21756 36642
rect 21700 36574 21756 36608
rect 21700 36540 21711 36574
rect 21745 36540 21756 36574
rect 21700 36506 21756 36540
rect 21700 36472 21711 36506
rect 21745 36472 21756 36506
rect 21700 36438 21756 36472
rect 21700 36404 21711 36438
rect 21745 36404 21756 36438
rect 21700 36370 21756 36404
rect 21700 36336 21711 36370
rect 21745 36336 21756 36370
rect 21700 36302 21756 36336
rect 21700 36268 21711 36302
rect 21745 36268 21756 36302
rect 21700 36234 21756 36268
rect 21700 36200 21711 36234
rect 21745 36200 21756 36234
rect 21700 36166 21756 36200
rect 21700 36132 21711 36166
rect 21745 36132 21756 36166
rect 21700 36098 21756 36132
rect 21700 36064 21711 36098
rect 21745 36064 21756 36098
rect 21700 36018 21756 36064
rect 22356 37322 22412 37368
rect 22356 37288 22367 37322
rect 22401 37288 22412 37322
rect 22356 37254 22412 37288
rect 22356 37220 22367 37254
rect 22401 37220 22412 37254
rect 22356 37186 22412 37220
rect 22356 37152 22367 37186
rect 22401 37152 22412 37186
rect 22356 37118 22412 37152
rect 22356 37084 22367 37118
rect 22401 37084 22412 37118
rect 22356 37050 22412 37084
rect 22356 37016 22367 37050
rect 22401 37016 22412 37050
rect 22356 36982 22412 37016
rect 22356 36948 22367 36982
rect 22401 36948 22412 36982
rect 22356 36914 22412 36948
rect 22356 36880 22367 36914
rect 22401 36880 22412 36914
rect 22356 36846 22412 36880
rect 22356 36812 22367 36846
rect 22401 36812 22412 36846
rect 22356 36778 22412 36812
rect 22356 36744 22367 36778
rect 22401 36744 22412 36778
rect 22356 36710 22412 36744
rect 22356 36676 22367 36710
rect 22401 36676 22412 36710
rect 22356 36642 22412 36676
rect 22356 36608 22367 36642
rect 22401 36608 22412 36642
rect 22356 36574 22412 36608
rect 22356 36540 22367 36574
rect 22401 36540 22412 36574
rect 22356 36506 22412 36540
rect 22356 36472 22367 36506
rect 22401 36472 22412 36506
rect 22356 36438 22412 36472
rect 22356 36404 22367 36438
rect 22401 36404 22412 36438
rect 22356 36370 22412 36404
rect 22356 36336 22367 36370
rect 22401 36336 22412 36370
rect 22356 36302 22412 36336
rect 22356 36268 22367 36302
rect 22401 36268 22412 36302
rect 22356 36234 22412 36268
rect 22356 36200 22367 36234
rect 22401 36200 22412 36234
rect 22356 36166 22412 36200
rect 22356 36132 22367 36166
rect 22401 36132 22412 36166
rect 22356 36098 22412 36132
rect 22356 36064 22367 36098
rect 22401 36064 22412 36098
rect 22356 36018 22412 36064
rect 23012 37322 23057 37368
rect 23012 37288 23023 37322
rect 23012 37254 23057 37288
rect 23012 37220 23023 37254
rect 23012 37186 23057 37220
rect 23012 37152 23023 37186
rect 23012 37118 23057 37152
rect 23012 37084 23023 37118
rect 23012 37050 23057 37084
rect 23012 37016 23023 37050
rect 23012 36982 23057 37016
rect 23012 36948 23023 36982
rect 23012 36914 23057 36948
rect 23012 36880 23023 36914
rect 23012 36846 23057 36880
rect 23012 36812 23023 36846
rect 23012 36778 23057 36812
rect 23012 36744 23023 36778
rect 23012 36710 23057 36744
rect 23012 36676 23023 36710
rect 23012 36642 23057 36676
rect 23012 36608 23023 36642
rect 23012 36574 23057 36608
rect 23012 36540 23023 36574
rect 23012 36506 23057 36540
rect 23012 36472 23023 36506
rect 23012 36438 23057 36472
rect 23012 36404 23023 36438
rect 23012 36370 23057 36404
rect 23012 36336 23023 36370
rect 23012 36302 23057 36336
rect 23012 36268 23023 36302
rect 23012 36234 23057 36268
rect 23012 36200 23023 36234
rect 23012 36166 23057 36200
rect 23012 36132 23023 36166
rect 23012 36098 23057 36132
rect 23012 36064 23023 36098
rect 23012 36018 23057 36064
rect 9767 34054 9820 34099
rect 9767 34020 9775 34054
rect 9809 34020 9820 34054
rect 9767 33986 9820 34020
rect 9767 33952 9775 33986
rect 9809 33952 9820 33986
rect 9767 33918 9820 33952
rect 9767 33884 9775 33918
rect 9809 33884 9820 33918
rect 9767 33850 9820 33884
rect 9767 33816 9775 33850
rect 9809 33816 9820 33850
rect 9767 33782 9820 33816
rect 9767 33748 9775 33782
rect 9809 33748 9820 33782
rect 9767 33714 9820 33748
rect 9767 33680 9775 33714
rect 9809 33680 9820 33714
rect 9767 33646 9820 33680
rect 9767 33612 9775 33646
rect 9809 33612 9820 33646
rect 9767 33578 9820 33612
rect 9767 33544 9775 33578
rect 9809 33544 9820 33578
rect 9767 33499 9820 33544
rect 10020 34054 10076 34099
rect 10020 34020 10031 34054
rect 10065 34020 10076 34054
rect 10020 33986 10076 34020
rect 10020 33952 10031 33986
rect 10065 33952 10076 33986
rect 10020 33918 10076 33952
rect 10020 33884 10031 33918
rect 10065 33884 10076 33918
rect 10020 33850 10076 33884
rect 10020 33816 10031 33850
rect 10065 33816 10076 33850
rect 10020 33782 10076 33816
rect 10020 33748 10031 33782
rect 10065 33748 10076 33782
rect 10020 33714 10076 33748
rect 10020 33680 10031 33714
rect 10065 33680 10076 33714
rect 10020 33646 10076 33680
rect 10020 33612 10031 33646
rect 10065 33612 10076 33646
rect 10020 33578 10076 33612
rect 10020 33544 10031 33578
rect 10065 33544 10076 33578
rect 10020 33499 10076 33544
rect 10276 34054 10332 34099
rect 10276 34020 10287 34054
rect 10321 34020 10332 34054
rect 10276 33986 10332 34020
rect 10276 33952 10287 33986
rect 10321 33952 10332 33986
rect 10276 33918 10332 33952
rect 10276 33884 10287 33918
rect 10321 33884 10332 33918
rect 10276 33850 10332 33884
rect 10276 33816 10287 33850
rect 10321 33816 10332 33850
rect 10276 33782 10332 33816
rect 10276 33748 10287 33782
rect 10321 33748 10332 33782
rect 10276 33714 10332 33748
rect 10276 33680 10287 33714
rect 10321 33680 10332 33714
rect 10276 33646 10332 33680
rect 10276 33612 10287 33646
rect 10321 33612 10332 33646
rect 10276 33578 10332 33612
rect 10276 33544 10287 33578
rect 10321 33544 10332 33578
rect 10276 33499 10332 33544
rect 10532 34054 10585 34099
rect 10532 34020 10543 34054
rect 10577 34020 10585 34054
rect 10532 33986 10585 34020
rect 10532 33952 10543 33986
rect 10577 33952 10585 33986
rect 10532 33918 10585 33952
rect 10532 33884 10543 33918
rect 10577 33884 10585 33918
rect 10532 33850 10585 33884
rect 10532 33816 10543 33850
rect 10577 33816 10585 33850
rect 10532 33782 10585 33816
rect 10532 33748 10543 33782
rect 10577 33748 10585 33782
rect 10532 33714 10585 33748
rect 10532 33680 10543 33714
rect 10577 33680 10585 33714
rect 10532 33646 10585 33680
rect 10532 33612 10543 33646
rect 10577 33612 10585 33646
rect 10532 33578 10585 33612
rect 10532 33544 10543 33578
rect 10577 33544 10585 33578
rect 10532 33499 10585 33544
rect 10641 34054 10694 34099
rect 10641 34020 10649 34054
rect 10683 34020 10694 34054
rect 10641 33986 10694 34020
rect 10641 33952 10649 33986
rect 10683 33952 10694 33986
rect 10641 33918 10694 33952
rect 10641 33884 10649 33918
rect 10683 33884 10694 33918
rect 10641 33850 10694 33884
rect 10641 33816 10649 33850
rect 10683 33816 10694 33850
rect 10641 33782 10694 33816
rect 10641 33748 10649 33782
rect 10683 33748 10694 33782
rect 10641 33714 10694 33748
rect 10641 33680 10649 33714
rect 10683 33680 10694 33714
rect 10641 33646 10694 33680
rect 10641 33612 10649 33646
rect 10683 33612 10694 33646
rect 10641 33578 10694 33612
rect 10641 33544 10649 33578
rect 10683 33544 10694 33578
rect 10641 33499 10694 33544
rect 10894 34054 10950 34099
rect 10894 34020 10905 34054
rect 10939 34020 10950 34054
rect 10894 33986 10950 34020
rect 10894 33952 10905 33986
rect 10939 33952 10950 33986
rect 10894 33918 10950 33952
rect 10894 33884 10905 33918
rect 10939 33884 10950 33918
rect 10894 33850 10950 33884
rect 10894 33816 10905 33850
rect 10939 33816 10950 33850
rect 10894 33782 10950 33816
rect 10894 33748 10905 33782
rect 10939 33748 10950 33782
rect 10894 33714 10950 33748
rect 10894 33680 10905 33714
rect 10939 33680 10950 33714
rect 10894 33646 10950 33680
rect 10894 33612 10905 33646
rect 10939 33612 10950 33646
rect 10894 33578 10950 33612
rect 10894 33544 10905 33578
rect 10939 33544 10950 33578
rect 10894 33499 10950 33544
rect 11150 34054 11206 34099
rect 11150 34020 11161 34054
rect 11195 34020 11206 34054
rect 11150 33986 11206 34020
rect 11150 33952 11161 33986
rect 11195 33952 11206 33986
rect 11150 33918 11206 33952
rect 11150 33884 11161 33918
rect 11195 33884 11206 33918
rect 11150 33850 11206 33884
rect 11150 33816 11161 33850
rect 11195 33816 11206 33850
rect 11150 33782 11206 33816
rect 11150 33748 11161 33782
rect 11195 33748 11206 33782
rect 11150 33714 11206 33748
rect 11150 33680 11161 33714
rect 11195 33680 11206 33714
rect 11150 33646 11206 33680
rect 11150 33612 11161 33646
rect 11195 33612 11206 33646
rect 11150 33578 11206 33612
rect 11150 33544 11161 33578
rect 11195 33544 11206 33578
rect 11150 33499 11206 33544
rect 11406 34054 11459 34099
rect 11406 34020 11417 34054
rect 11451 34020 11459 34054
rect 11406 33986 11459 34020
rect 11406 33952 11417 33986
rect 11451 33952 11459 33986
rect 11406 33918 11459 33952
rect 11406 33884 11417 33918
rect 11451 33884 11459 33918
rect 11406 33850 11459 33884
rect 11406 33816 11417 33850
rect 11451 33816 11459 33850
rect 11406 33782 11459 33816
rect 11406 33748 11417 33782
rect 11451 33748 11459 33782
rect 11406 33714 11459 33748
rect 11406 33680 11417 33714
rect 11451 33680 11459 33714
rect 11406 33646 11459 33680
rect 11406 33612 11417 33646
rect 11451 33612 11459 33646
rect 11406 33578 11459 33612
rect 11406 33544 11417 33578
rect 11451 33544 11459 33578
rect 11406 33499 11459 33544
rect 11955 34092 12008 34124
rect 11955 34058 11963 34092
rect 11997 34058 12008 34092
rect 11955 34024 12008 34058
rect 11955 33990 11963 34024
rect 11997 33990 12008 34024
rect 11955 33956 12008 33990
rect 11955 33922 11963 33956
rect 11997 33922 12008 33956
rect 11955 33888 12008 33922
rect 11955 33854 11963 33888
rect 11997 33854 12008 33888
rect 11955 33820 12008 33854
rect 11955 33786 11963 33820
rect 11997 33786 12008 33820
rect 11955 33752 12008 33786
rect 11955 33718 11963 33752
rect 11997 33718 12008 33752
rect 11955 33684 12008 33718
rect 11955 33650 11963 33684
rect 11997 33650 12008 33684
rect 11955 33616 12008 33650
rect 11955 33582 11963 33616
rect 11997 33582 12008 33616
rect 11955 33548 12008 33582
rect 11955 33514 11963 33548
rect 11997 33514 12008 33548
rect 11955 33480 12008 33514
rect 11955 33446 11963 33480
rect 11997 33446 12008 33480
rect 11955 33414 12008 33446
rect 12208 34092 12264 34124
rect 12208 34058 12219 34092
rect 12253 34058 12264 34092
rect 12208 34024 12264 34058
rect 12208 33990 12219 34024
rect 12253 33990 12264 34024
rect 12208 33956 12264 33990
rect 12208 33922 12219 33956
rect 12253 33922 12264 33956
rect 12208 33888 12264 33922
rect 12208 33854 12219 33888
rect 12253 33854 12264 33888
rect 12208 33820 12264 33854
rect 12208 33786 12219 33820
rect 12253 33786 12264 33820
rect 12208 33752 12264 33786
rect 12208 33718 12219 33752
rect 12253 33718 12264 33752
rect 12208 33684 12264 33718
rect 12208 33650 12219 33684
rect 12253 33650 12264 33684
rect 12208 33616 12264 33650
rect 12208 33582 12219 33616
rect 12253 33582 12264 33616
rect 12208 33548 12264 33582
rect 12208 33514 12219 33548
rect 12253 33514 12264 33548
rect 12208 33480 12264 33514
rect 12208 33446 12219 33480
rect 12253 33446 12264 33480
rect 12208 33414 12264 33446
rect 12464 34092 12520 34124
rect 12464 34058 12475 34092
rect 12509 34058 12520 34092
rect 12464 34024 12520 34058
rect 12464 33990 12475 34024
rect 12509 33990 12520 34024
rect 12464 33956 12520 33990
rect 12464 33922 12475 33956
rect 12509 33922 12520 33956
rect 12464 33888 12520 33922
rect 12464 33854 12475 33888
rect 12509 33854 12520 33888
rect 12464 33820 12520 33854
rect 12464 33786 12475 33820
rect 12509 33786 12520 33820
rect 12464 33752 12520 33786
rect 12464 33718 12475 33752
rect 12509 33718 12520 33752
rect 12464 33684 12520 33718
rect 12464 33650 12475 33684
rect 12509 33650 12520 33684
rect 12464 33616 12520 33650
rect 12464 33582 12475 33616
rect 12509 33582 12520 33616
rect 12464 33548 12520 33582
rect 12464 33514 12475 33548
rect 12509 33514 12520 33548
rect 12464 33480 12520 33514
rect 12464 33446 12475 33480
rect 12509 33446 12520 33480
rect 12464 33414 12520 33446
rect 12720 34092 12773 34124
rect 12720 34058 12731 34092
rect 12765 34058 12773 34092
rect 12720 34024 12773 34058
rect 12720 33990 12731 34024
rect 12765 33990 12773 34024
rect 12720 33956 12773 33990
rect 12720 33922 12731 33956
rect 12765 33922 12773 33956
rect 12720 33888 12773 33922
rect 12720 33854 12731 33888
rect 12765 33854 12773 33888
rect 12720 33820 12773 33854
rect 12720 33786 12731 33820
rect 12765 33786 12773 33820
rect 12720 33752 12773 33786
rect 12720 33718 12731 33752
rect 12765 33718 12773 33752
rect 12720 33684 12773 33718
rect 12720 33650 12731 33684
rect 12765 33650 12773 33684
rect 12720 33616 12773 33650
rect 12720 33582 12731 33616
rect 12765 33582 12773 33616
rect 12720 33548 12773 33582
rect 12720 33514 12731 33548
rect 12765 33514 12773 33548
rect 12720 33480 12773 33514
rect 12720 33446 12731 33480
rect 12765 33446 12773 33480
rect 12720 33414 12773 33446
rect 13089 34057 13142 34106
rect 13089 34023 13097 34057
rect 13131 34023 13142 34057
rect 13089 33989 13142 34023
rect 13089 33955 13097 33989
rect 13131 33955 13142 33989
rect 13089 33921 13142 33955
rect 13089 33887 13097 33921
rect 13131 33887 13142 33921
rect 13089 33853 13142 33887
rect 13089 33819 13097 33853
rect 13131 33819 13142 33853
rect 13089 33785 13142 33819
rect 13089 33751 13097 33785
rect 13131 33751 13142 33785
rect 13089 33717 13142 33751
rect 13089 33683 13097 33717
rect 13131 33683 13142 33717
rect 13089 33649 13142 33683
rect 13089 33615 13097 33649
rect 13131 33615 13142 33649
rect 13089 33581 13142 33615
rect 13089 33547 13097 33581
rect 13131 33547 13142 33581
rect 13089 33513 13142 33547
rect 13089 33479 13097 33513
rect 13131 33479 13142 33513
rect 13089 33431 13142 33479
rect 13742 34057 13795 34106
rect 13742 34023 13753 34057
rect 13787 34023 13795 34057
rect 13742 33989 13795 34023
rect 13742 33955 13753 33989
rect 13787 33955 13795 33989
rect 13742 33921 13795 33955
rect 13742 33887 13753 33921
rect 13787 33887 13795 33921
rect 13742 33853 13795 33887
rect 13742 33819 13753 33853
rect 13787 33819 13795 33853
rect 13742 33785 13795 33819
rect 13742 33751 13753 33785
rect 13787 33751 13795 33785
rect 13742 33717 13795 33751
rect 13742 33683 13753 33717
rect 13787 33683 13795 33717
rect 13742 33649 13795 33683
rect 13742 33615 13753 33649
rect 13787 33615 13795 33649
rect 13742 33581 13795 33615
rect 13742 33547 13753 33581
rect 13787 33547 13795 33581
rect 13742 33513 13795 33547
rect 13742 33479 13753 33513
rect 13787 33479 13795 33513
rect 13742 33431 13795 33479
rect 13867 34057 13920 34106
rect 13867 34023 13875 34057
rect 13909 34023 13920 34057
rect 13867 33989 13920 34023
rect 13867 33955 13875 33989
rect 13909 33955 13920 33989
rect 13867 33921 13920 33955
rect 13867 33887 13875 33921
rect 13909 33887 13920 33921
rect 13867 33853 13920 33887
rect 13867 33819 13875 33853
rect 13909 33819 13920 33853
rect 13867 33785 13920 33819
rect 13867 33751 13875 33785
rect 13909 33751 13920 33785
rect 13867 33717 13920 33751
rect 13867 33683 13875 33717
rect 13909 33683 13920 33717
rect 13867 33649 13920 33683
rect 13867 33615 13875 33649
rect 13909 33615 13920 33649
rect 13867 33581 13920 33615
rect 13867 33547 13875 33581
rect 13909 33547 13920 33581
rect 13867 33513 13920 33547
rect 13867 33479 13875 33513
rect 13909 33479 13920 33513
rect 13867 33431 13920 33479
rect 14520 34057 14565 34106
rect 14520 34023 14531 34057
rect 14520 33989 14565 34023
rect 14520 33955 14531 33989
rect 14520 33921 14565 33955
rect 14520 33887 14531 33921
rect 14520 33853 14565 33887
rect 14520 33819 14531 33853
rect 14520 33785 14565 33819
rect 14520 33751 14531 33785
rect 14520 33717 14565 33751
rect 14520 33683 14531 33717
rect 14520 33649 14565 33683
rect 14520 33615 14531 33649
rect 14520 33581 14565 33615
rect 14520 33547 14531 33581
rect 14520 33513 14565 33547
rect 14520 33479 14531 33513
rect 14520 33431 14565 33479
<< ndiffc >>
rect 9629 32723 9663 32757
rect 9629 32655 9663 32689
rect 9629 32587 9663 32621
rect 9629 32519 9663 32553
rect 9629 32451 9663 32485
rect 9629 32383 9663 32417
rect 9629 32315 9663 32349
rect 9629 32247 9663 32281
rect 9629 32179 9663 32213
rect 9629 32111 9663 32145
rect 9629 32043 9663 32077
rect 9629 31975 9663 32009
rect 9629 31907 9663 31941
rect 9629 31839 9663 31873
rect 9629 31771 9663 31805
rect 9629 31703 9663 31737
rect 9629 31635 9663 31669
rect 9629 31567 9663 31601
rect 9629 31499 9663 31533
rect 9629 31431 9663 31465
rect 9985 32723 10019 32757
rect 9985 32655 10019 32689
rect 9985 32587 10019 32621
rect 9985 32519 10019 32553
rect 9985 32451 10019 32485
rect 9985 32383 10019 32417
rect 9985 32315 10019 32349
rect 9985 32247 10019 32281
rect 9985 32179 10019 32213
rect 9985 32111 10019 32145
rect 9985 32043 10019 32077
rect 9985 31975 10019 32009
rect 9985 31907 10019 31941
rect 9985 31839 10019 31873
rect 9985 31771 10019 31805
rect 9985 31703 10019 31737
rect 9985 31635 10019 31669
rect 9985 31567 10019 31601
rect 9985 31499 10019 31533
rect 9985 31431 10019 31465
rect 10341 32723 10375 32757
rect 10341 32655 10375 32689
rect 10341 32587 10375 32621
rect 10341 32519 10375 32553
rect 10341 32451 10375 32485
rect 10341 32383 10375 32417
rect 10341 32315 10375 32349
rect 10341 32247 10375 32281
rect 10341 32179 10375 32213
rect 10341 32111 10375 32145
rect 10341 32043 10375 32077
rect 10341 31975 10375 32009
rect 10341 31907 10375 31941
rect 10341 31839 10375 31873
rect 10341 31771 10375 31805
rect 10341 31703 10375 31737
rect 10341 31635 10375 31669
rect 10341 31567 10375 31601
rect 10341 31499 10375 31533
rect 10341 31431 10375 31465
rect 10697 32723 10731 32757
rect 10697 32655 10731 32689
rect 10697 32587 10731 32621
rect 10697 32519 10731 32553
rect 10697 32451 10731 32485
rect 10697 32383 10731 32417
rect 10697 32315 10731 32349
rect 10697 32247 10731 32281
rect 10697 32179 10731 32213
rect 10697 32111 10731 32145
rect 10697 32043 10731 32077
rect 10697 31975 10731 32009
rect 10697 31907 10731 31941
rect 10697 31839 10731 31873
rect 10697 31771 10731 31805
rect 10697 31703 10731 31737
rect 10697 31635 10731 31669
rect 10697 31567 10731 31601
rect 10697 31499 10731 31533
rect 10697 31431 10731 31465
rect 11053 32723 11087 32757
rect 11053 32655 11087 32689
rect 11053 32587 11087 32621
rect 11053 32519 11087 32553
rect 11053 32451 11087 32485
rect 11053 32383 11087 32417
rect 11053 32315 11087 32349
rect 11053 32247 11087 32281
rect 11053 32179 11087 32213
rect 11053 32111 11087 32145
rect 11053 32043 11087 32077
rect 11053 31975 11087 32009
rect 11053 31907 11087 31941
rect 11053 31839 11087 31873
rect 11053 31771 11087 31805
rect 11053 31703 11087 31737
rect 11053 31635 11087 31669
rect 11053 31567 11087 31601
rect 11053 31499 11087 31533
rect 11053 31431 11087 31465
rect 11450 32785 11484 32819
rect 11450 32717 11484 32751
rect 11450 32649 11484 32683
rect 11450 32581 11484 32615
rect 11450 32513 11484 32547
rect 11450 32445 11484 32479
rect 11450 32377 11484 32411
rect 12006 32785 12040 32819
rect 12006 32717 12040 32751
rect 12006 32649 12040 32683
rect 12006 32581 12040 32615
rect 12006 32513 12040 32547
rect 12006 32445 12040 32479
rect 12006 32377 12040 32411
rect 12562 32785 12596 32819
rect 12562 32717 12596 32751
rect 12562 32649 12596 32683
rect 12562 32581 12596 32615
rect 12562 32513 12596 32547
rect 12562 32445 12596 32479
rect 12562 32377 12596 32411
rect 13118 32785 13152 32819
rect 13118 32717 13152 32751
rect 13118 32649 13152 32683
rect 13118 32581 13152 32615
rect 13118 32513 13152 32547
rect 13118 32445 13152 32479
rect 13118 32377 13152 32411
rect 13224 32785 13258 32819
rect 13224 32717 13258 32751
rect 13224 32649 13258 32683
rect 13224 32581 13258 32615
rect 13224 32513 13258 32547
rect 13224 32445 13258 32479
rect 13224 32377 13258 32411
rect 13780 32785 13814 32819
rect 13780 32717 13814 32751
rect 13780 32649 13814 32683
rect 13780 32581 13814 32615
rect 13780 32513 13814 32547
rect 13780 32445 13814 32479
rect 13780 32377 13814 32411
rect 14336 32785 14370 32819
rect 14336 32717 14370 32751
rect 14336 32649 14370 32683
rect 14336 32581 14370 32615
rect 14336 32513 14370 32547
rect 14336 32445 14370 32479
rect 14336 32377 14370 32411
rect 11450 32231 11484 32265
rect 11450 32163 11484 32197
rect 11450 32095 11484 32129
rect 11450 32027 11484 32061
rect 11450 31959 11484 31993
rect 11450 31891 11484 31925
rect 11450 31823 11484 31857
rect 12006 32231 12040 32265
rect 12006 32163 12040 32197
rect 12006 32095 12040 32129
rect 12006 32027 12040 32061
rect 12006 31959 12040 31993
rect 12006 31891 12040 31925
rect 12006 31823 12040 31857
rect 12562 32231 12596 32265
rect 12562 32163 12596 32197
rect 12562 32095 12596 32129
rect 12562 32027 12596 32061
rect 12562 31959 12596 31993
rect 12562 31891 12596 31925
rect 12562 31823 12596 31857
rect 13118 32231 13152 32265
rect 13118 32163 13152 32197
rect 13118 32095 13152 32129
rect 13118 32027 13152 32061
rect 13118 31959 13152 31993
rect 13118 31891 13152 31925
rect 13118 31823 13152 31857
rect 13224 32231 13258 32265
rect 13224 32163 13258 32197
rect 13224 32095 13258 32129
rect 13224 32027 13258 32061
rect 13224 31959 13258 31993
rect 13224 31891 13258 31925
rect 13224 31823 13258 31857
rect 13780 32231 13814 32265
rect 13780 32163 13814 32197
rect 13780 32095 13814 32129
rect 13780 32027 13814 32061
rect 13780 31959 13814 31993
rect 13780 31891 13814 31925
rect 13780 31823 13814 31857
rect 14336 32231 14370 32265
rect 14336 32163 14370 32197
rect 14336 32095 14370 32129
rect 14336 32027 14370 32061
rect 14336 31959 14370 31993
rect 14336 31891 14370 31925
rect 14336 31823 14370 31857
rect 9629 31009 9663 31043
rect 9629 30941 9663 30975
rect 9629 30873 9663 30907
rect 9629 30805 9663 30839
rect 9629 30737 9663 30771
rect 9629 30669 9663 30703
rect 9629 30601 9663 30635
rect 9629 30533 9663 30567
rect 9629 30465 9663 30499
rect 9629 30397 9663 30431
rect 9629 30329 9663 30363
rect 9629 30261 9663 30295
rect 9629 30193 9663 30227
rect 9629 30125 9663 30159
rect 9629 30057 9663 30091
rect 9629 29989 9663 30023
rect 9629 29921 9663 29955
rect 9629 29853 9663 29887
rect 9629 29785 9663 29819
rect 9629 29717 9663 29751
rect 9985 31009 10019 31043
rect 9985 30941 10019 30975
rect 9985 30873 10019 30907
rect 9985 30805 10019 30839
rect 9985 30737 10019 30771
rect 9985 30669 10019 30703
rect 9985 30601 10019 30635
rect 9985 30533 10019 30567
rect 9985 30465 10019 30499
rect 9985 30397 10019 30431
rect 9985 30329 10019 30363
rect 9985 30261 10019 30295
rect 9985 30193 10019 30227
rect 9985 30125 10019 30159
rect 9985 30057 10019 30091
rect 9985 29989 10019 30023
rect 9985 29921 10019 29955
rect 9985 29853 10019 29887
rect 9985 29785 10019 29819
rect 9985 29717 10019 29751
rect 10341 31009 10375 31043
rect 10341 30941 10375 30975
rect 10341 30873 10375 30907
rect 10341 30805 10375 30839
rect 10341 30737 10375 30771
rect 10341 30669 10375 30703
rect 10341 30601 10375 30635
rect 10341 30533 10375 30567
rect 10341 30465 10375 30499
rect 10341 30397 10375 30431
rect 10341 30329 10375 30363
rect 10341 30261 10375 30295
rect 10341 30193 10375 30227
rect 10341 30125 10375 30159
rect 10341 30057 10375 30091
rect 10341 29989 10375 30023
rect 10341 29921 10375 29955
rect 10341 29853 10375 29887
rect 10341 29785 10375 29819
rect 10341 29717 10375 29751
rect 10697 31009 10731 31043
rect 10697 30941 10731 30975
rect 10697 30873 10731 30907
rect 10697 30805 10731 30839
rect 10697 30737 10731 30771
rect 10697 30669 10731 30703
rect 10697 30601 10731 30635
rect 10697 30533 10731 30567
rect 10697 30465 10731 30499
rect 10697 30397 10731 30431
rect 10697 30329 10731 30363
rect 10697 30261 10731 30295
rect 10697 30193 10731 30227
rect 10697 30125 10731 30159
rect 10697 30057 10731 30091
rect 10697 29989 10731 30023
rect 10697 29921 10731 29955
rect 10697 29853 10731 29887
rect 10697 29785 10731 29819
rect 10697 29717 10731 29751
rect 11053 31009 11087 31043
rect 11053 30941 11087 30975
rect 11053 30873 11087 30907
rect 11053 30805 11087 30839
rect 11053 30737 11087 30771
rect 11053 30669 11087 30703
rect 11053 30601 11087 30635
rect 11053 30533 11087 30567
rect 11053 30465 11087 30499
rect 11053 30397 11087 30431
rect 11053 30329 11087 30363
rect 11053 30261 11087 30295
rect 11053 30193 11087 30227
rect 11053 30125 11087 30159
rect 11053 30057 11087 30091
rect 11053 29989 11087 30023
rect 11053 29921 11087 29955
rect 11053 29853 11087 29887
rect 11053 29785 11087 29819
rect 11053 29717 11087 29751
<< pdiffc >>
rect 9577 37306 9611 37340
rect 9577 37238 9611 37272
rect 9577 37170 9611 37204
rect 9577 37102 9611 37136
rect 9577 37034 9611 37068
rect 9577 36966 9611 37000
rect 9577 36898 9611 36932
rect 9577 36830 9611 36864
rect 9577 36762 9611 36796
rect 9577 36694 9611 36728
rect 9577 36626 9611 36660
rect 9577 36558 9611 36592
rect 9577 36490 9611 36524
rect 9577 36422 9611 36456
rect 9577 36354 9611 36388
rect 9577 36286 9611 36320
rect 9577 36218 9611 36252
rect 9577 36150 9611 36184
rect 9577 36082 9611 36116
rect 10233 37306 10267 37340
rect 10233 37238 10267 37272
rect 10233 37170 10267 37204
rect 10233 37102 10267 37136
rect 10233 37034 10267 37068
rect 10233 36966 10267 37000
rect 10233 36898 10267 36932
rect 10233 36830 10267 36864
rect 10233 36762 10267 36796
rect 10233 36694 10267 36728
rect 10233 36626 10267 36660
rect 10233 36558 10267 36592
rect 10233 36490 10267 36524
rect 10233 36422 10267 36456
rect 10233 36354 10267 36388
rect 10233 36286 10267 36320
rect 10233 36218 10267 36252
rect 10233 36150 10267 36184
rect 10233 36082 10267 36116
rect 10339 37306 10373 37340
rect 10339 37238 10373 37272
rect 10339 37170 10373 37204
rect 10339 37102 10373 37136
rect 10339 37034 10373 37068
rect 10339 36966 10373 37000
rect 10339 36898 10373 36932
rect 10339 36830 10373 36864
rect 10339 36762 10373 36796
rect 10339 36694 10373 36728
rect 10339 36626 10373 36660
rect 10339 36558 10373 36592
rect 10339 36490 10373 36524
rect 10339 36422 10373 36456
rect 10339 36354 10373 36388
rect 10339 36286 10373 36320
rect 10339 36218 10373 36252
rect 10339 36150 10373 36184
rect 10339 36082 10373 36116
rect 10995 37306 11029 37340
rect 10995 37238 11029 37272
rect 10995 37170 11029 37204
rect 10995 37102 11029 37136
rect 10995 37034 11029 37068
rect 10995 36966 11029 37000
rect 10995 36898 11029 36932
rect 10995 36830 11029 36864
rect 10995 36762 11029 36796
rect 10995 36694 11029 36728
rect 10995 36626 11029 36660
rect 10995 36558 11029 36592
rect 10995 36490 11029 36524
rect 10995 36422 11029 36456
rect 10995 36354 11029 36388
rect 10995 36286 11029 36320
rect 10995 36218 11029 36252
rect 10995 36150 11029 36184
rect 10995 36082 11029 36116
rect 11651 37306 11685 37340
rect 11651 37238 11685 37272
rect 11651 37170 11685 37204
rect 11651 37102 11685 37136
rect 11651 37034 11685 37068
rect 11651 36966 11685 37000
rect 11651 36898 11685 36932
rect 11651 36830 11685 36864
rect 11651 36762 11685 36796
rect 11651 36694 11685 36728
rect 11651 36626 11685 36660
rect 11651 36558 11685 36592
rect 11651 36490 11685 36524
rect 11651 36422 11685 36456
rect 11651 36354 11685 36388
rect 11651 36286 11685 36320
rect 11651 36218 11685 36252
rect 11651 36150 11685 36184
rect 11651 36082 11685 36116
rect 12307 37306 12341 37340
rect 12307 37238 12341 37272
rect 12307 37170 12341 37204
rect 12307 37102 12341 37136
rect 12307 37034 12341 37068
rect 12307 36966 12341 37000
rect 12307 36898 12341 36932
rect 12307 36830 12341 36864
rect 12307 36762 12341 36796
rect 12307 36694 12341 36728
rect 12307 36626 12341 36660
rect 12307 36558 12341 36592
rect 12307 36490 12341 36524
rect 12307 36422 12341 36456
rect 12307 36354 12341 36388
rect 12307 36286 12341 36320
rect 12307 36218 12341 36252
rect 12307 36150 12341 36184
rect 12307 36082 12341 36116
rect 12963 37306 12997 37340
rect 12963 37238 12997 37272
rect 12963 37170 12997 37204
rect 12963 37102 12997 37136
rect 12963 37034 12997 37068
rect 12963 36966 12997 37000
rect 12963 36898 12997 36932
rect 12963 36830 12997 36864
rect 12963 36762 12997 36796
rect 12963 36694 12997 36728
rect 12963 36626 12997 36660
rect 12963 36558 12997 36592
rect 12963 36490 12997 36524
rect 12963 36422 12997 36456
rect 12963 36354 12997 36388
rect 12963 36286 12997 36320
rect 12963 36218 12997 36252
rect 12963 36150 12997 36184
rect 12963 36082 12997 36116
rect 13619 37306 13653 37340
rect 13619 37238 13653 37272
rect 13619 37170 13653 37204
rect 13619 37102 13653 37136
rect 13619 37034 13653 37068
rect 13619 36966 13653 37000
rect 13619 36898 13653 36932
rect 13619 36830 13653 36864
rect 13619 36762 13653 36796
rect 13619 36694 13653 36728
rect 13619 36626 13653 36660
rect 13619 36558 13653 36592
rect 13619 36490 13653 36524
rect 13619 36422 13653 36456
rect 13619 36354 13653 36388
rect 13619 36286 13653 36320
rect 13619 36218 13653 36252
rect 13619 36150 13653 36184
rect 13619 36082 13653 36116
rect 14275 37306 14309 37340
rect 14275 37238 14309 37272
rect 14275 37170 14309 37204
rect 14275 37102 14309 37136
rect 14275 37034 14309 37068
rect 14275 36966 14309 37000
rect 14275 36898 14309 36932
rect 14275 36830 14309 36864
rect 14275 36762 14309 36796
rect 14275 36694 14309 36728
rect 14275 36626 14309 36660
rect 14275 36558 14309 36592
rect 14275 36490 14309 36524
rect 14275 36422 14309 36456
rect 14275 36354 14309 36388
rect 14275 36286 14309 36320
rect 14275 36218 14309 36252
rect 14275 36150 14309 36184
rect 14275 36082 14309 36116
rect 9577 35884 9611 35918
rect 9577 35816 9611 35850
rect 9577 35748 9611 35782
rect 9577 35680 9611 35714
rect 9577 35612 9611 35646
rect 9577 35544 9611 35578
rect 9577 35476 9611 35510
rect 9577 35408 9611 35442
rect 9577 35340 9611 35374
rect 9577 35272 9611 35306
rect 9577 35204 9611 35238
rect 9577 35136 9611 35170
rect 9577 35068 9611 35102
rect 9577 35000 9611 35034
rect 9577 34932 9611 34966
rect 9577 34864 9611 34898
rect 9577 34796 9611 34830
rect 9577 34728 9611 34762
rect 9577 34660 9611 34694
rect 10233 35884 10267 35918
rect 10233 35816 10267 35850
rect 10233 35748 10267 35782
rect 10233 35680 10267 35714
rect 10233 35612 10267 35646
rect 10233 35544 10267 35578
rect 10233 35476 10267 35510
rect 10233 35408 10267 35442
rect 10233 35340 10267 35374
rect 10233 35272 10267 35306
rect 10233 35204 10267 35238
rect 10233 35136 10267 35170
rect 10233 35068 10267 35102
rect 10233 35000 10267 35034
rect 10233 34932 10267 34966
rect 10233 34864 10267 34898
rect 10233 34796 10267 34830
rect 10233 34728 10267 34762
rect 10233 34660 10267 34694
rect 10339 35884 10373 35918
rect 10339 35816 10373 35850
rect 10339 35748 10373 35782
rect 10339 35680 10373 35714
rect 10339 35612 10373 35646
rect 10339 35544 10373 35578
rect 10339 35476 10373 35510
rect 10339 35408 10373 35442
rect 10339 35340 10373 35374
rect 10339 35272 10373 35306
rect 10339 35204 10373 35238
rect 10339 35136 10373 35170
rect 10339 35068 10373 35102
rect 10339 35000 10373 35034
rect 10339 34932 10373 34966
rect 10339 34864 10373 34898
rect 10339 34796 10373 34830
rect 10339 34728 10373 34762
rect 10339 34660 10373 34694
rect 10995 35884 11029 35918
rect 10995 35816 11029 35850
rect 10995 35748 11029 35782
rect 10995 35680 11029 35714
rect 10995 35612 11029 35646
rect 10995 35544 11029 35578
rect 10995 35476 11029 35510
rect 10995 35408 11029 35442
rect 10995 35340 11029 35374
rect 10995 35272 11029 35306
rect 10995 35204 11029 35238
rect 10995 35136 11029 35170
rect 10995 35068 11029 35102
rect 10995 35000 11029 35034
rect 10995 34932 11029 34966
rect 10995 34864 11029 34898
rect 10995 34796 11029 34830
rect 10995 34728 11029 34762
rect 10995 34660 11029 34694
rect 11651 35884 11685 35918
rect 11651 35816 11685 35850
rect 11651 35748 11685 35782
rect 11651 35680 11685 35714
rect 11651 35612 11685 35646
rect 11651 35544 11685 35578
rect 11651 35476 11685 35510
rect 11651 35408 11685 35442
rect 11651 35340 11685 35374
rect 11651 35272 11685 35306
rect 11651 35204 11685 35238
rect 11651 35136 11685 35170
rect 11651 35068 11685 35102
rect 11651 35000 11685 35034
rect 11651 34932 11685 34966
rect 11651 34864 11685 34898
rect 11651 34796 11685 34830
rect 11651 34728 11685 34762
rect 11651 34660 11685 34694
rect 12307 35884 12341 35918
rect 12307 35816 12341 35850
rect 12307 35748 12341 35782
rect 12307 35680 12341 35714
rect 12307 35612 12341 35646
rect 12307 35544 12341 35578
rect 12307 35476 12341 35510
rect 12307 35408 12341 35442
rect 12307 35340 12341 35374
rect 12307 35272 12341 35306
rect 12307 35204 12341 35238
rect 12307 35136 12341 35170
rect 12307 35068 12341 35102
rect 12307 35000 12341 35034
rect 12307 34932 12341 34966
rect 12307 34864 12341 34898
rect 12307 34796 12341 34830
rect 12307 34728 12341 34762
rect 12307 34660 12341 34694
rect 12963 35884 12997 35918
rect 12963 35816 12997 35850
rect 12963 35748 12997 35782
rect 12963 35680 12997 35714
rect 12963 35612 12997 35646
rect 12963 35544 12997 35578
rect 12963 35476 12997 35510
rect 12963 35408 12997 35442
rect 12963 35340 12997 35374
rect 12963 35272 12997 35306
rect 12963 35204 12997 35238
rect 12963 35136 12997 35170
rect 12963 35068 12997 35102
rect 12963 35000 12997 35034
rect 12963 34932 12997 34966
rect 12963 34864 12997 34898
rect 12963 34796 12997 34830
rect 12963 34728 12997 34762
rect 12963 34660 12997 34694
rect 13619 35884 13653 35918
rect 13619 35816 13653 35850
rect 13619 35748 13653 35782
rect 13619 35680 13653 35714
rect 13619 35612 13653 35646
rect 13619 35544 13653 35578
rect 13619 35476 13653 35510
rect 13619 35408 13653 35442
rect 13619 35340 13653 35374
rect 13619 35272 13653 35306
rect 13619 35204 13653 35238
rect 13619 35136 13653 35170
rect 13619 35068 13653 35102
rect 13619 35000 13653 35034
rect 13619 34932 13653 34966
rect 13619 34864 13653 34898
rect 13619 34796 13653 34830
rect 13619 34728 13653 34762
rect 13619 34660 13653 34694
rect 14275 35884 14309 35918
rect 14275 35816 14309 35850
rect 14275 35748 14309 35782
rect 14275 35680 14309 35714
rect 14275 35612 14309 35646
rect 14275 35544 14309 35578
rect 14275 35476 14309 35510
rect 14275 35408 14309 35442
rect 14275 35340 14309 35374
rect 14275 35272 14309 35306
rect 14275 35204 14309 35238
rect 14275 35136 14309 35170
rect 14275 35068 14309 35102
rect 14275 35000 14309 35034
rect 14275 34932 14309 34966
rect 14275 34864 14309 34898
rect 14275 34796 14309 34830
rect 14275 34728 14309 34762
rect 14275 34660 14309 34694
rect 19087 37288 19121 37322
rect 19087 37220 19121 37254
rect 19087 37152 19121 37186
rect 19087 37084 19121 37118
rect 19087 37016 19121 37050
rect 19087 36948 19121 36982
rect 19087 36880 19121 36914
rect 19087 36812 19121 36846
rect 19087 36744 19121 36778
rect 19087 36676 19121 36710
rect 19087 36608 19121 36642
rect 19087 36540 19121 36574
rect 19087 36472 19121 36506
rect 19087 36404 19121 36438
rect 19087 36336 19121 36370
rect 19087 36268 19121 36302
rect 19087 36200 19121 36234
rect 19087 36132 19121 36166
rect 19087 36064 19121 36098
rect 19743 37288 19777 37322
rect 19743 37220 19777 37254
rect 19743 37152 19777 37186
rect 19743 37084 19777 37118
rect 19743 37016 19777 37050
rect 19743 36948 19777 36982
rect 19743 36880 19777 36914
rect 19743 36812 19777 36846
rect 19743 36744 19777 36778
rect 19743 36676 19777 36710
rect 19743 36608 19777 36642
rect 19743 36540 19777 36574
rect 19743 36472 19777 36506
rect 19743 36404 19777 36438
rect 19743 36336 19777 36370
rect 19743 36268 19777 36302
rect 19743 36200 19777 36234
rect 19743 36132 19777 36166
rect 19743 36064 19777 36098
rect 20399 37288 20433 37322
rect 20399 37220 20433 37254
rect 20399 37152 20433 37186
rect 20399 37084 20433 37118
rect 20399 37016 20433 37050
rect 20399 36948 20433 36982
rect 20399 36880 20433 36914
rect 20399 36812 20433 36846
rect 20399 36744 20433 36778
rect 20399 36676 20433 36710
rect 20399 36608 20433 36642
rect 20399 36540 20433 36574
rect 20399 36472 20433 36506
rect 20399 36404 20433 36438
rect 20399 36336 20433 36370
rect 20399 36268 20433 36302
rect 20399 36200 20433 36234
rect 20399 36132 20433 36166
rect 20399 36064 20433 36098
rect 21055 37288 21089 37322
rect 21055 37220 21089 37254
rect 21055 37152 21089 37186
rect 21055 37084 21089 37118
rect 21055 37016 21089 37050
rect 21055 36948 21089 36982
rect 21055 36880 21089 36914
rect 21055 36812 21089 36846
rect 21055 36744 21089 36778
rect 21055 36676 21089 36710
rect 21055 36608 21089 36642
rect 21055 36540 21089 36574
rect 21055 36472 21089 36506
rect 21055 36404 21089 36438
rect 21055 36336 21089 36370
rect 21055 36268 21089 36302
rect 21055 36200 21089 36234
rect 21055 36132 21089 36166
rect 21055 36064 21089 36098
rect 21711 37288 21745 37322
rect 21711 37220 21745 37254
rect 21711 37152 21745 37186
rect 21711 37084 21745 37118
rect 21711 37016 21745 37050
rect 21711 36948 21745 36982
rect 21711 36880 21745 36914
rect 21711 36812 21745 36846
rect 21711 36744 21745 36778
rect 21711 36676 21745 36710
rect 21711 36608 21745 36642
rect 21711 36540 21745 36574
rect 21711 36472 21745 36506
rect 21711 36404 21745 36438
rect 21711 36336 21745 36370
rect 21711 36268 21745 36302
rect 21711 36200 21745 36234
rect 21711 36132 21745 36166
rect 21711 36064 21745 36098
rect 22367 37288 22401 37322
rect 22367 37220 22401 37254
rect 22367 37152 22401 37186
rect 22367 37084 22401 37118
rect 22367 37016 22401 37050
rect 22367 36948 22401 36982
rect 22367 36880 22401 36914
rect 22367 36812 22401 36846
rect 22367 36744 22401 36778
rect 22367 36676 22401 36710
rect 22367 36608 22401 36642
rect 22367 36540 22401 36574
rect 22367 36472 22401 36506
rect 22367 36404 22401 36438
rect 22367 36336 22401 36370
rect 22367 36268 22401 36302
rect 22367 36200 22401 36234
rect 22367 36132 22401 36166
rect 22367 36064 22401 36098
rect 23023 37288 23057 37322
rect 23023 37220 23057 37254
rect 23023 37152 23057 37186
rect 23023 37084 23057 37118
rect 23023 37016 23057 37050
rect 23023 36948 23057 36982
rect 23023 36880 23057 36914
rect 23023 36812 23057 36846
rect 23023 36744 23057 36778
rect 23023 36676 23057 36710
rect 23023 36608 23057 36642
rect 23023 36540 23057 36574
rect 23023 36472 23057 36506
rect 23023 36404 23057 36438
rect 23023 36336 23057 36370
rect 23023 36268 23057 36302
rect 23023 36200 23057 36234
rect 23023 36132 23057 36166
rect 23023 36064 23057 36098
rect 9775 34020 9809 34054
rect 9775 33952 9809 33986
rect 9775 33884 9809 33918
rect 9775 33816 9809 33850
rect 9775 33748 9809 33782
rect 9775 33680 9809 33714
rect 9775 33612 9809 33646
rect 9775 33544 9809 33578
rect 10031 34020 10065 34054
rect 10031 33952 10065 33986
rect 10031 33884 10065 33918
rect 10031 33816 10065 33850
rect 10031 33748 10065 33782
rect 10031 33680 10065 33714
rect 10031 33612 10065 33646
rect 10031 33544 10065 33578
rect 10287 34020 10321 34054
rect 10287 33952 10321 33986
rect 10287 33884 10321 33918
rect 10287 33816 10321 33850
rect 10287 33748 10321 33782
rect 10287 33680 10321 33714
rect 10287 33612 10321 33646
rect 10287 33544 10321 33578
rect 10543 34020 10577 34054
rect 10543 33952 10577 33986
rect 10543 33884 10577 33918
rect 10543 33816 10577 33850
rect 10543 33748 10577 33782
rect 10543 33680 10577 33714
rect 10543 33612 10577 33646
rect 10543 33544 10577 33578
rect 10649 34020 10683 34054
rect 10649 33952 10683 33986
rect 10649 33884 10683 33918
rect 10649 33816 10683 33850
rect 10649 33748 10683 33782
rect 10649 33680 10683 33714
rect 10649 33612 10683 33646
rect 10649 33544 10683 33578
rect 10905 34020 10939 34054
rect 10905 33952 10939 33986
rect 10905 33884 10939 33918
rect 10905 33816 10939 33850
rect 10905 33748 10939 33782
rect 10905 33680 10939 33714
rect 10905 33612 10939 33646
rect 10905 33544 10939 33578
rect 11161 34020 11195 34054
rect 11161 33952 11195 33986
rect 11161 33884 11195 33918
rect 11161 33816 11195 33850
rect 11161 33748 11195 33782
rect 11161 33680 11195 33714
rect 11161 33612 11195 33646
rect 11161 33544 11195 33578
rect 11417 34020 11451 34054
rect 11417 33952 11451 33986
rect 11417 33884 11451 33918
rect 11417 33816 11451 33850
rect 11417 33748 11451 33782
rect 11417 33680 11451 33714
rect 11417 33612 11451 33646
rect 11417 33544 11451 33578
rect 11963 34058 11997 34092
rect 11963 33990 11997 34024
rect 11963 33922 11997 33956
rect 11963 33854 11997 33888
rect 11963 33786 11997 33820
rect 11963 33718 11997 33752
rect 11963 33650 11997 33684
rect 11963 33582 11997 33616
rect 11963 33514 11997 33548
rect 11963 33446 11997 33480
rect 12219 34058 12253 34092
rect 12219 33990 12253 34024
rect 12219 33922 12253 33956
rect 12219 33854 12253 33888
rect 12219 33786 12253 33820
rect 12219 33718 12253 33752
rect 12219 33650 12253 33684
rect 12219 33582 12253 33616
rect 12219 33514 12253 33548
rect 12219 33446 12253 33480
rect 12475 34058 12509 34092
rect 12475 33990 12509 34024
rect 12475 33922 12509 33956
rect 12475 33854 12509 33888
rect 12475 33786 12509 33820
rect 12475 33718 12509 33752
rect 12475 33650 12509 33684
rect 12475 33582 12509 33616
rect 12475 33514 12509 33548
rect 12475 33446 12509 33480
rect 12731 34058 12765 34092
rect 12731 33990 12765 34024
rect 12731 33922 12765 33956
rect 12731 33854 12765 33888
rect 12731 33786 12765 33820
rect 12731 33718 12765 33752
rect 12731 33650 12765 33684
rect 12731 33582 12765 33616
rect 12731 33514 12765 33548
rect 12731 33446 12765 33480
rect 13097 34023 13131 34057
rect 13097 33955 13131 33989
rect 13097 33887 13131 33921
rect 13097 33819 13131 33853
rect 13097 33751 13131 33785
rect 13097 33683 13131 33717
rect 13097 33615 13131 33649
rect 13097 33547 13131 33581
rect 13097 33479 13131 33513
rect 13753 34023 13787 34057
rect 13753 33955 13787 33989
rect 13753 33887 13787 33921
rect 13753 33819 13787 33853
rect 13753 33751 13787 33785
rect 13753 33683 13787 33717
rect 13753 33615 13787 33649
rect 13753 33547 13787 33581
rect 13753 33479 13787 33513
rect 13875 34023 13909 34057
rect 13875 33955 13909 33989
rect 13875 33887 13909 33921
rect 13875 33819 13909 33853
rect 13875 33751 13909 33785
rect 13875 33683 13909 33717
rect 13875 33615 13909 33649
rect 13875 33547 13909 33581
rect 13875 33479 13909 33513
rect 14531 34023 14565 34057
rect 14531 33955 14565 33989
rect 14531 33887 14565 33921
rect 14531 33819 14565 33853
rect 14531 33751 14565 33785
rect 14531 33683 14565 33717
rect 14531 33615 14565 33649
rect 14531 33547 14565 33581
rect 14531 33479 14565 33513
<< psubdiff >>
rect 7638 33092 7662 33098
rect 6952 33058 6976 33092
rect 7010 33058 7044 33092
rect 7078 33058 7112 33092
rect 7146 33058 7180 33092
rect 7214 33058 7248 33092
rect 7282 33058 7316 33092
rect 7350 33058 7384 33092
rect 7418 33058 7452 33092
rect 7486 33058 7520 33092
rect 7554 33064 7662 33092
rect 7696 33064 7730 33098
rect 7764 33064 7798 33098
rect 7832 33092 7924 33098
rect 7832 33064 7914 33092
rect 7554 33058 7672 33064
rect 7890 33058 7914 33064
rect 7948 33058 8036 33092
rect 6952 32976 6986 33058
rect 8002 33040 8036 33058
rect 6952 32908 6986 32942
rect 8002 33016 8072 33040
rect 8002 33006 8038 33016
rect 8038 32948 8072 32982
rect 6952 32840 6986 32874
rect 6952 32772 6986 32806
rect 6952 32704 6986 32738
rect 6952 32636 6986 32670
rect 6952 32568 6986 32602
rect 6952 32500 6986 32534
rect 6952 32432 6986 32466
rect 6952 32364 6986 32398
rect 6952 32296 6986 32330
rect 6952 32228 6986 32262
rect 6952 32160 6986 32194
rect 6952 32092 6986 32126
rect 6952 32024 6986 32058
rect 6952 31956 6986 31990
rect 6854 31898 6878 31932
rect 6912 31922 6952 31932
rect 6912 31898 6986 31922
rect 8038 32880 8072 32914
rect 9434 33004 9458 33038
rect 9492 33004 9526 33038
rect 9560 33004 9594 33038
rect 9628 33004 9662 33038
rect 9696 33004 9730 33038
rect 9764 33004 9798 33038
rect 9832 33004 9866 33038
rect 9900 33004 9934 33038
rect 9968 33004 10002 33038
rect 10036 33004 10070 33038
rect 10104 33004 10138 33038
rect 10172 33004 10206 33038
rect 10240 33004 10274 33038
rect 10308 33004 10342 33038
rect 10376 33004 10410 33038
rect 10444 33004 10478 33038
rect 10512 33004 10546 33038
rect 10580 33004 10614 33038
rect 10648 33004 10682 33038
rect 10716 33004 10750 33038
rect 10784 33004 10818 33038
rect 10852 33004 10886 33038
rect 10920 33004 10954 33038
rect 10988 33004 11022 33038
rect 11056 33004 11090 33038
rect 11124 33004 11158 33038
rect 11192 33014 11276 33038
rect 11192 33004 11242 33014
rect 9434 32927 9468 33004
rect 11242 32946 11276 32980
rect 8038 32812 8072 32846
rect 8038 32744 8072 32778
rect 9434 32859 9468 32893
rect 9621 32910 11095 32922
rect 9621 32876 9650 32910
rect 9684 32876 9718 32910
rect 9752 32876 9786 32910
rect 9820 32876 9854 32910
rect 9888 32876 9922 32910
rect 9956 32876 10044 32910
rect 10078 32876 10112 32910
rect 10146 32876 10180 32910
rect 10214 32876 10248 32910
rect 10282 32876 10400 32910
rect 10434 32876 10468 32910
rect 10502 32876 10536 32910
rect 10570 32876 10604 32910
rect 10638 32876 10743 32910
rect 10777 32876 10811 32910
rect 10845 32876 10879 32910
rect 10913 32876 10947 32910
rect 10981 32876 11015 32910
rect 11049 32876 11095 32910
rect 9621 32864 11095 32876
rect 11242 32878 11276 32912
rect 9434 32791 9468 32825
rect 11242 32810 11276 32844
rect 8038 32676 8072 32710
rect 9434 32723 9468 32757
rect 8038 32608 8072 32642
rect 8038 32540 8072 32574
rect 8038 32472 8072 32506
rect 8038 32404 8072 32438
rect 8038 32336 8072 32370
rect 8038 32268 8072 32302
rect 8038 32200 8072 32234
rect 8038 32132 8072 32166
rect 8038 32064 8072 32098
rect 8038 31963 8072 32030
rect 6854 31827 6888 31898
rect 6854 31759 6888 31793
rect 6854 31691 6888 31725
rect 6854 31623 6888 31657
rect 8038 31895 8072 31929
rect 8038 31827 8072 31861
rect 8038 31759 8072 31793
rect 8038 31691 8072 31725
rect 8038 31623 8072 31657
rect 6888 31589 6928 31599
rect 6854 31565 6928 31589
rect 6962 31565 6996 31599
rect 7030 31565 7064 31599
rect 7098 31565 7132 31599
rect 7166 31565 7200 31599
rect 7234 31565 7268 31599
rect 7302 31565 7336 31599
rect 7370 31565 7394 31599
rect 7360 31468 7394 31565
rect 7360 31400 7394 31434
rect 7360 31332 7394 31366
rect 7360 31264 7394 31298
rect 7360 31196 7394 31230
rect 7360 31128 7394 31162
rect 7360 31060 7394 31094
rect 7360 30992 7394 31026
rect 7331 30958 7360 30968
rect 7331 30934 7394 30958
rect 8038 31555 8072 31589
rect 8038 31487 8072 31521
rect 8038 31419 8072 31453
rect 8038 31351 8072 31385
rect 8038 31283 8072 31317
rect 8038 31215 8072 31249
rect 8038 31147 8072 31181
rect 8038 31079 8072 31113
rect 8038 30968 8072 31045
rect 9434 32655 9468 32689
rect 9434 32587 9468 32621
rect 9434 32519 9468 32553
rect 9434 32451 9468 32485
rect 9434 32383 9468 32417
rect 9434 32315 9468 32349
rect 9434 32247 9468 32281
rect 9434 32179 9468 32213
rect 9434 32111 9468 32145
rect 9434 32043 9468 32077
rect 9434 31975 9468 32009
rect 9434 31907 9468 31941
rect 9434 31839 9468 31873
rect 9434 31771 9468 31805
rect 9434 31703 9468 31737
rect 9434 31635 9468 31669
rect 9434 31567 9468 31601
rect 9434 31499 9468 31533
rect 9434 31431 9468 31465
rect 9434 31363 9468 31397
rect 11242 32742 11276 32776
rect 11242 32674 11276 32708
rect 11242 32606 11276 32640
rect 11242 32538 11276 32572
rect 11242 32470 11276 32504
rect 11242 32402 11276 32436
rect 11242 32334 11276 32368
rect 11242 32266 11276 32300
rect 11242 32198 11276 32232
rect 11242 32130 11276 32164
rect 11242 32062 11276 32096
rect 11242 31994 11276 32028
rect 11242 31926 11276 31960
rect 11242 31858 11276 31892
rect 11242 31790 11276 31824
rect 11242 31722 11276 31756
rect 11242 31654 11276 31688
rect 11242 31586 11276 31620
rect 11330 33014 11422 33038
rect 11364 33004 11422 33014
rect 11456 33004 11490 33038
rect 11524 33004 11558 33038
rect 11592 33004 11626 33038
rect 11660 33004 11694 33038
rect 11728 33004 11762 33038
rect 11796 33004 11830 33038
rect 11864 33004 11898 33038
rect 11932 33004 11966 33038
rect 12000 33004 12034 33038
rect 12068 33004 12102 33038
rect 12136 33004 12170 33038
rect 12204 33004 12238 33038
rect 12272 33004 12306 33038
rect 12340 33004 12374 33038
rect 12408 33004 12442 33038
rect 12476 33004 12510 33038
rect 12544 33004 12578 33038
rect 12612 33004 12646 33038
rect 12680 33004 12714 33038
rect 12748 33004 12782 33038
rect 12816 33004 12850 33038
rect 12884 33004 12918 33038
rect 12952 33004 12986 33038
rect 13020 33004 13054 33038
rect 13088 33004 13122 33038
rect 13156 33004 13190 33038
rect 13224 33004 13258 33038
rect 13292 33004 13326 33038
rect 13360 33004 13394 33038
rect 13428 33004 13462 33038
rect 13496 33004 13530 33038
rect 13564 33004 13598 33038
rect 13632 33004 13666 33038
rect 13700 33004 13734 33038
rect 13768 33004 13802 33038
rect 13836 33004 13870 33038
rect 13904 33004 13938 33038
rect 13972 33004 14006 33038
rect 14040 33004 14074 33038
rect 14108 33004 14142 33038
rect 14176 33004 14210 33038
rect 14244 33004 14278 33038
rect 14312 33004 14346 33038
rect 14380 33004 14414 33038
rect 14448 33004 14482 33038
rect 14516 33004 14550 33038
rect 14584 33004 14618 33038
rect 14652 33004 14686 33038
rect 14720 33004 14754 33038
rect 14788 33004 14822 33038
rect 14856 33004 14890 33038
rect 14924 33004 14958 33038
rect 14992 33004 15026 33038
rect 15060 33004 15094 33038
rect 15128 33004 15162 33038
rect 15196 33004 15230 33038
rect 15264 33004 15298 33038
rect 15332 33004 15366 33038
rect 15400 33004 15434 33038
rect 15468 33004 15502 33038
rect 15536 33004 15570 33038
rect 15604 33004 15638 33038
rect 15672 33004 15706 33038
rect 15740 33004 15774 33038
rect 15808 33004 15842 33038
rect 15876 33004 15910 33038
rect 15944 33004 15978 33038
rect 16012 33004 16046 33038
rect 16080 33004 16114 33038
rect 16148 33004 16182 33038
rect 16216 33004 16250 33038
rect 16284 33004 16318 33038
rect 16352 33004 16376 33038
rect 11330 32946 11364 32980
rect 16342 32970 16376 33004
rect 11330 32878 11364 32912
rect 16342 32902 16376 32936
rect 11330 32810 11364 32844
rect 11330 32742 11364 32776
rect 11330 32674 11364 32708
rect 11330 32606 11364 32640
rect 11330 32538 11364 32572
rect 11330 32470 11364 32504
rect 11330 32402 11364 32436
rect 11330 32334 11364 32368
rect 16342 32834 16376 32868
rect 16342 32766 16376 32800
rect 16342 32698 16376 32732
rect 16342 32630 16376 32664
rect 16342 32562 16376 32596
rect 16342 32494 16376 32528
rect 16342 32426 16376 32460
rect 16342 32358 16376 32392
rect 11330 32266 11364 32300
rect 11330 32198 11364 32232
rect 11330 32130 11364 32164
rect 11330 32062 11364 32096
rect 11330 31994 11364 32028
rect 11330 31926 11364 31960
rect 11330 31858 11364 31892
rect 11330 31790 11364 31824
rect 16342 32290 16376 32324
rect 16342 32222 16376 32256
rect 16342 32154 16376 32188
rect 16342 32086 16376 32120
rect 16342 32018 16376 32052
rect 16342 31950 16376 31984
rect 16342 31882 16376 31916
rect 16342 31814 16376 31848
rect 11330 31722 11364 31756
rect 16342 31746 16376 31780
rect 11330 31654 11364 31688
rect 11442 31712 13160 31724
rect 11442 31678 11469 31712
rect 11503 31678 11537 31712
rect 11571 31678 11605 31712
rect 11639 31678 11673 31712
rect 11707 31678 11741 31712
rect 11775 31678 11809 31712
rect 11843 31678 11877 31712
rect 11911 31678 11945 31712
rect 11979 31678 12063 31712
rect 12097 31678 12131 31712
rect 12165 31678 12199 31712
rect 12233 31678 12267 31712
rect 12301 31678 12335 31712
rect 12369 31678 12403 31712
rect 12437 31678 12471 31712
rect 12505 31678 12606 31712
rect 12640 31678 12674 31712
rect 12708 31678 12742 31712
rect 12776 31678 12810 31712
rect 12844 31678 12878 31712
rect 12912 31678 12946 31712
rect 12980 31678 13014 31712
rect 13048 31678 13082 31712
rect 13116 31678 13160 31712
rect 11442 31666 13160 31678
rect 13216 31712 14378 31724
rect 13216 31678 13260 31712
rect 13294 31678 13328 31712
rect 13362 31678 13396 31712
rect 13430 31678 13464 31712
rect 13498 31678 13532 31712
rect 13566 31678 13600 31712
rect 13634 31678 13668 31712
rect 13702 31678 13736 31712
rect 13770 31678 13841 31712
rect 13875 31678 13909 31712
rect 13943 31678 13977 31712
rect 14011 31678 14045 31712
rect 14079 31678 14113 31712
rect 14147 31678 14181 31712
rect 14215 31678 14249 31712
rect 14283 31678 14317 31712
rect 14351 31678 14378 31712
rect 13216 31666 14378 31678
rect 16342 31678 16376 31712
rect 11330 31586 11364 31620
rect 16342 31610 16376 31644
rect 11330 31552 11354 31586
rect 11388 31552 11422 31586
rect 11456 31552 11490 31586
rect 11524 31552 11558 31586
rect 11592 31552 11626 31586
rect 11660 31552 11694 31586
rect 11728 31552 11762 31586
rect 11796 31552 11830 31586
rect 11864 31552 11898 31586
rect 11932 31552 11966 31586
rect 12000 31552 12034 31586
rect 12068 31552 12102 31586
rect 12136 31552 12170 31586
rect 12204 31552 12238 31586
rect 12272 31552 12306 31586
rect 12340 31552 12374 31586
rect 12408 31552 12442 31586
rect 12476 31552 12510 31586
rect 12544 31552 12578 31586
rect 12612 31552 12646 31586
rect 12680 31552 12714 31586
rect 12748 31552 12782 31586
rect 12816 31552 12850 31586
rect 12884 31552 12918 31586
rect 12952 31552 12986 31586
rect 13020 31552 13054 31586
rect 13088 31552 13122 31586
rect 13156 31552 13190 31586
rect 13224 31552 13258 31586
rect 13292 31552 13326 31586
rect 13360 31552 13394 31586
rect 13428 31552 13462 31586
rect 13496 31552 13530 31586
rect 13564 31552 13598 31586
rect 13632 31552 13666 31586
rect 13700 31552 13734 31586
rect 13768 31552 13877 31586
rect 13911 31552 13945 31586
rect 13979 31552 14013 31586
rect 14047 31552 14081 31586
rect 14115 31552 14149 31586
rect 14183 31552 14217 31586
rect 14251 31552 14285 31586
rect 14319 31552 14353 31586
rect 14387 31552 14421 31586
rect 14455 31552 14489 31586
rect 14523 31552 14557 31586
rect 14591 31552 14625 31586
rect 14659 31552 14693 31586
rect 14727 31552 14761 31586
rect 14795 31552 14829 31586
rect 14863 31552 14897 31586
rect 14931 31552 14965 31586
rect 14999 31552 15033 31586
rect 15067 31552 15101 31586
rect 15135 31552 15169 31586
rect 15203 31552 15237 31586
rect 15271 31552 15305 31586
rect 15339 31552 15373 31586
rect 15407 31552 15441 31586
rect 15475 31552 15509 31586
rect 15543 31552 15577 31586
rect 15611 31552 15645 31586
rect 15679 31552 15713 31586
rect 15747 31552 15781 31586
rect 15815 31552 15849 31586
rect 15883 31552 15917 31586
rect 15951 31552 15985 31586
rect 16019 31552 16053 31586
rect 16087 31552 16121 31586
rect 16155 31552 16189 31586
rect 16223 31552 16257 31586
rect 16291 31576 16342 31586
rect 16291 31552 16376 31576
rect 11242 31518 11276 31552
rect 11242 31450 11276 31484
rect 9434 31295 9468 31329
rect 11242 31382 11276 31416
rect 11242 31314 11276 31348
rect 9434 31194 9468 31261
rect 11242 31246 11276 31280
rect 11242 31178 11276 31212
rect 12668 31346 12777 31380
rect 12811 31346 12845 31380
rect 12879 31346 12913 31380
rect 12947 31346 12981 31380
rect 13015 31346 13049 31380
rect 13083 31346 13117 31380
rect 13151 31346 13185 31380
rect 13219 31346 13253 31380
rect 13287 31346 13321 31380
rect 13355 31346 13389 31380
rect 13423 31346 13457 31380
rect 13491 31346 13525 31380
rect 13559 31346 13593 31380
rect 13627 31346 13661 31380
rect 13695 31346 13729 31380
rect 13763 31346 13797 31380
rect 13831 31346 13865 31380
rect 13899 31346 13933 31380
rect 13967 31346 14001 31380
rect 14035 31346 14069 31380
rect 14103 31346 14137 31380
rect 14171 31346 14205 31380
rect 14239 31346 14273 31380
rect 14307 31346 14341 31380
rect 14375 31346 14409 31380
rect 14443 31346 14477 31380
rect 14511 31346 14620 31380
rect 12668 31266 12702 31346
rect 14586 31266 14620 31346
rect 9434 31126 9468 31160
rect 9434 31058 9468 31092
rect 11242 31110 11276 31144
rect 12668 31198 12702 31232
rect 14586 31198 14620 31232
rect 9434 30990 9468 31024
rect 8038 30944 8101 30968
rect 8038 30934 8067 30944
rect 7331 30843 7365 30934
rect 7331 30775 7365 30809
rect 7331 30707 7365 30741
rect 8067 30876 8101 30910
rect 8067 30808 8101 30842
rect 8067 30683 8101 30774
rect 7365 30673 7431 30683
rect 7331 30649 7431 30673
rect 7465 30649 7499 30683
rect 7533 30649 7567 30683
rect 7601 30649 7635 30683
rect 7669 30649 7703 30683
rect 7737 30649 7771 30683
rect 7805 30649 7839 30683
rect 7873 30649 7907 30683
rect 7941 30649 7975 30683
rect 8009 30649 8043 30683
rect 8077 30649 8101 30683
rect 9434 30922 9468 30956
rect 9434 30854 9468 30888
rect 9434 30786 9468 30820
rect 9434 30718 9468 30752
rect 9434 30650 9468 30684
rect 9434 30582 9468 30616
rect 9434 30514 9468 30548
rect 9434 30446 9468 30480
rect 9434 30378 9468 30412
rect 9434 30310 9468 30344
rect 9434 30242 9468 30276
rect 9434 30174 9468 30208
rect 9434 30106 9468 30140
rect 9434 30038 9468 30072
rect 9434 29970 9468 30004
rect 9434 29902 9468 29936
rect 9434 29834 9468 29868
rect 9434 29766 9468 29800
rect 9434 29698 9468 29732
rect 11242 31042 11276 31076
rect 12668 31084 12702 31164
rect 14586 31084 14620 31164
rect 12668 31050 12777 31084
rect 12811 31050 12845 31084
rect 12879 31050 12913 31084
rect 12947 31050 12981 31084
rect 13015 31050 13049 31084
rect 13083 31050 13117 31084
rect 13151 31050 13185 31084
rect 13219 31050 13253 31084
rect 13287 31050 13321 31084
rect 13355 31050 13389 31084
rect 13423 31050 13457 31084
rect 13491 31050 13525 31084
rect 13559 31050 13593 31084
rect 13627 31050 13661 31084
rect 13695 31050 13729 31084
rect 13763 31050 13797 31084
rect 13831 31050 13865 31084
rect 13899 31050 13933 31084
rect 13967 31050 14001 31084
rect 14035 31050 14069 31084
rect 14103 31050 14137 31084
rect 14171 31050 14205 31084
rect 14239 31050 14273 31084
rect 14307 31050 14341 31084
rect 14375 31050 14409 31084
rect 14443 31050 14477 31084
rect 14511 31050 14620 31084
rect 11242 30974 11276 31008
rect 11242 30906 11276 30940
rect 11242 30838 11276 30872
rect 11242 30770 11276 30804
rect 11242 30702 11276 30736
rect 11242 30634 11276 30668
rect 11242 30566 11276 30600
rect 11242 30498 11276 30532
rect 11242 30430 11276 30464
rect 11242 30362 11276 30396
rect 11242 30294 11276 30328
rect 11242 30226 11276 30260
rect 11242 30158 11276 30192
rect 11242 30090 11276 30124
rect 11242 30022 11276 30056
rect 11242 29954 11276 29988
rect 11242 29886 11276 29920
rect 11242 29818 11276 29852
rect 11242 29750 11276 29784
rect 11242 29682 11276 29716
rect 9434 29630 9468 29664
rect 11242 29614 11276 29648
rect 9434 29562 9468 29596
rect 9621 29598 11095 29610
rect 9621 29564 9667 29598
rect 9701 29564 9735 29598
rect 9769 29564 9803 29598
rect 9837 29564 9871 29598
rect 9905 29564 9939 29598
rect 9973 29564 10078 29598
rect 10112 29564 10146 29598
rect 10180 29564 10214 29598
rect 10248 29564 10282 29598
rect 10316 29564 10417 29598
rect 10451 29564 10485 29598
rect 10519 29564 10553 29598
rect 10587 29564 10621 29598
rect 10655 29564 10743 29598
rect 10777 29564 10811 29598
rect 10845 29564 10879 29598
rect 10913 29564 10947 29598
rect 10981 29564 11015 29598
rect 11049 29564 11095 29598
rect 9621 29552 11095 29564
rect 9434 29494 9468 29528
rect 11242 29546 11276 29580
rect 11242 29470 11276 29512
rect 9468 29460 9518 29470
rect 9434 29436 9518 29460
rect 9552 29436 9586 29470
rect 9620 29436 9654 29470
rect 9688 29436 9722 29470
rect 9756 29436 9790 29470
rect 9824 29436 9858 29470
rect 9892 29436 9926 29470
rect 9960 29436 9994 29470
rect 10028 29436 10062 29470
rect 10096 29436 10130 29470
rect 10164 29436 10198 29470
rect 10232 29436 10266 29470
rect 10300 29436 10334 29470
rect 10368 29436 10402 29470
rect 10436 29436 10470 29470
rect 10504 29436 10538 29470
rect 10572 29436 10606 29470
rect 10640 29436 10674 29470
rect 10708 29436 10742 29470
rect 10776 29436 10810 29470
rect 10844 29436 10878 29470
rect 10912 29436 10946 29470
rect 10980 29436 11014 29470
rect 11048 29436 11082 29470
rect 11116 29436 11150 29470
rect 11184 29436 11218 29470
rect 11252 29436 11276 29470
rect 9650 14716 9674 14722
rect 8964 14682 8988 14716
rect 9022 14682 9056 14716
rect 9090 14682 9124 14716
rect 9158 14682 9192 14716
rect 9226 14682 9260 14716
rect 9294 14682 9328 14716
rect 9362 14682 9396 14716
rect 9430 14682 9464 14716
rect 9498 14682 9532 14716
rect 9566 14688 9674 14716
rect 9708 14688 9742 14722
rect 9776 14688 9810 14722
rect 9844 14716 9936 14722
rect 9844 14688 9926 14716
rect 9566 14682 9684 14688
rect 9902 14682 9926 14688
rect 9960 14682 10048 14716
rect 8964 14600 8998 14682
rect 10014 14664 10048 14682
rect 8964 14532 8998 14566
rect 10014 14640 10084 14664
rect 10014 14630 10050 14640
rect 10050 14572 10084 14606
rect 8964 14464 8998 14498
rect 8964 14396 8998 14430
rect 8964 14328 8998 14362
rect 8964 14260 8998 14294
rect 8964 14192 8998 14226
rect 8964 14124 8998 14158
rect 8964 14056 8998 14090
rect 8964 13988 8998 14022
rect 8964 13920 8998 13954
rect 8964 13852 8998 13886
rect 8964 13784 8998 13818
rect 8964 13716 8998 13750
rect 8964 13648 8998 13682
rect 8964 13580 8998 13614
rect 8866 13522 8890 13556
rect 8924 13546 8964 13556
rect 8924 13522 8998 13546
rect 10050 14504 10084 14538
rect 11446 14628 11470 14662
rect 11504 14628 11538 14662
rect 11572 14628 11606 14662
rect 11640 14628 11674 14662
rect 11708 14628 11742 14662
rect 11776 14628 11810 14662
rect 11844 14628 11878 14662
rect 11912 14628 11946 14662
rect 11980 14628 12014 14662
rect 12048 14628 12082 14662
rect 12116 14628 12150 14662
rect 12184 14628 12218 14662
rect 12252 14628 12286 14662
rect 12320 14628 12354 14662
rect 12388 14628 12422 14662
rect 12456 14628 12490 14662
rect 12524 14628 12558 14662
rect 12592 14628 12626 14662
rect 12660 14628 12694 14662
rect 12728 14628 12762 14662
rect 12796 14628 12830 14662
rect 12864 14628 12898 14662
rect 12932 14628 12966 14662
rect 13000 14628 13034 14662
rect 13068 14628 13102 14662
rect 13136 14628 13170 14662
rect 13204 14638 13288 14662
rect 13204 14628 13254 14638
rect 11446 14551 11480 14628
rect 10050 14436 10084 14470
rect 10050 14368 10084 14402
rect 11446 14483 11480 14517
rect 11446 14415 11480 14449
rect 10050 14300 10084 14334
rect 11446 14347 11480 14381
rect 10050 14232 10084 14266
rect 10050 14164 10084 14198
rect 10050 14096 10084 14130
rect 10050 14028 10084 14062
rect 10050 13960 10084 13994
rect 10050 13892 10084 13926
rect 10050 13824 10084 13858
rect 10050 13756 10084 13790
rect 10050 13688 10084 13722
rect 10050 13587 10084 13654
rect 8866 13451 8900 13522
rect 8866 13383 8900 13417
rect 8866 13315 8900 13349
rect 8866 13247 8900 13281
rect 10050 13519 10084 13553
rect 10050 13451 10084 13485
rect 10050 13383 10084 13417
rect 10050 13315 10084 13349
rect 10050 13247 10084 13281
rect 8900 13213 8940 13223
rect 8866 13189 8940 13213
rect 8974 13189 9008 13223
rect 9042 13189 9076 13223
rect 9110 13189 9144 13223
rect 9178 13189 9212 13223
rect 9246 13189 9280 13223
rect 9314 13189 9348 13223
rect 9382 13189 9406 13223
rect 9372 13092 9406 13189
rect 9372 13024 9406 13058
rect 9372 12956 9406 12990
rect 9372 12888 9406 12922
rect 9372 12820 9406 12854
rect 9372 12752 9406 12786
rect 9372 12684 9406 12718
rect 9372 12616 9406 12650
rect 9343 12582 9372 12592
rect 9343 12558 9406 12582
rect 10050 13179 10084 13213
rect 10050 13111 10084 13145
rect 10050 13043 10084 13077
rect 10050 12975 10084 13009
rect 10050 12907 10084 12941
rect 10050 12839 10084 12873
rect 10050 12771 10084 12805
rect 10050 12703 10084 12737
rect 10050 12592 10084 12669
rect 11446 14279 11480 14313
rect 11446 14211 11480 14245
rect 11446 14143 11480 14177
rect 11446 14075 11480 14109
rect 11446 14007 11480 14041
rect 11446 13939 11480 13973
rect 11446 13871 11480 13905
rect 11446 13803 11480 13837
rect 11446 13735 11480 13769
rect 11446 13667 11480 13701
rect 11446 13599 11480 13633
rect 11446 13531 11480 13565
rect 11446 13463 11480 13497
rect 11446 13395 11480 13429
rect 11446 13327 11480 13361
rect 11446 13259 11480 13293
rect 11446 13191 11480 13225
rect 11446 13123 11480 13157
rect 11446 13055 11480 13089
rect 11446 12987 11480 13021
rect 11446 12919 11480 12953
rect 11446 12818 11480 12885
rect 11446 12750 11480 12784
rect 11446 12682 11480 12716
rect 11446 12614 11480 12648
rect 10050 12568 10113 12592
rect 10050 12558 10079 12568
rect 9343 12467 9377 12558
rect 9343 12399 9377 12433
rect 9343 12331 9377 12365
rect 10079 12500 10113 12534
rect 10079 12432 10113 12466
rect 10079 12307 10113 12398
rect 9377 12297 9443 12307
rect 9343 12273 9443 12297
rect 9477 12273 9511 12307
rect 9545 12273 9579 12307
rect 9613 12273 9647 12307
rect 9681 12273 9715 12307
rect 9749 12273 9783 12307
rect 9817 12273 9851 12307
rect 9885 12273 9919 12307
rect 9953 12273 9987 12307
rect 10021 12273 10055 12307
rect 10089 12273 10113 12307
rect 11446 12546 11480 12580
rect 11446 12478 11480 12512
rect 11446 12410 11480 12444
rect 11446 12342 11480 12376
rect 11446 12274 11480 12308
rect 11446 12206 11480 12240
rect 11446 12138 11480 12172
rect 11446 12070 11480 12104
rect 11446 12002 11480 12036
rect 11446 11934 11480 11968
rect 11446 11866 11480 11900
rect 11446 11798 11480 11832
rect 11446 11730 11480 11764
rect 11446 11662 11480 11696
rect 11446 11594 11480 11628
rect 11446 11526 11480 11560
rect 11446 11458 11480 11492
rect 11446 11390 11480 11424
rect 11446 11322 11480 11356
rect 11446 11254 11480 11288
rect 11446 11186 11480 11220
rect 11446 11118 11480 11152
rect 13254 14570 13288 14604
rect 13254 14502 13288 14536
rect 13254 14434 13288 14468
rect 13254 14366 13288 14400
rect 13254 14298 13288 14332
rect 13254 14230 13288 14264
rect 13254 14162 13288 14196
rect 13254 14094 13288 14128
rect 13254 14026 13288 14060
rect 13254 13958 13288 13992
rect 13254 13890 13288 13924
rect 13254 13822 13288 13856
rect 13254 13754 13288 13788
rect 13254 13686 13288 13720
rect 13254 13618 13288 13652
rect 13254 13550 13288 13584
rect 13254 13482 13288 13516
rect 13254 13414 13288 13448
rect 13254 13346 13288 13380
rect 13254 13278 13288 13312
rect 13254 13210 13288 13244
rect 13342 14638 13434 14662
rect 13376 14628 13434 14638
rect 13468 14628 13502 14662
rect 13536 14628 13570 14662
rect 13604 14628 13638 14662
rect 13672 14628 13706 14662
rect 13740 14628 13774 14662
rect 13808 14628 13842 14662
rect 13876 14628 13910 14662
rect 13944 14628 13978 14662
rect 14012 14628 14046 14662
rect 14080 14628 14114 14662
rect 14148 14628 14182 14662
rect 14216 14628 14250 14662
rect 14284 14628 14318 14662
rect 14352 14628 14386 14662
rect 14420 14628 14454 14662
rect 14488 14628 14522 14662
rect 14556 14628 14590 14662
rect 14624 14628 14658 14662
rect 14692 14628 14726 14662
rect 14760 14628 14794 14662
rect 14828 14628 14862 14662
rect 14896 14628 14930 14662
rect 14964 14628 14998 14662
rect 15032 14628 15066 14662
rect 15100 14628 15134 14662
rect 15168 14628 15202 14662
rect 15236 14628 15270 14662
rect 15304 14628 15338 14662
rect 15372 14628 15406 14662
rect 15440 14628 15474 14662
rect 15508 14628 15542 14662
rect 15576 14628 15610 14662
rect 15644 14628 15678 14662
rect 15712 14628 15746 14662
rect 15780 14628 15814 14662
rect 15848 14628 15882 14662
rect 15916 14628 15950 14662
rect 15984 14628 16018 14662
rect 16052 14628 16086 14662
rect 16120 14628 16154 14662
rect 16188 14628 16222 14662
rect 16256 14628 16290 14662
rect 16324 14628 16358 14662
rect 16392 14628 16426 14662
rect 16460 14628 16494 14662
rect 16528 14628 16562 14662
rect 16596 14628 16630 14662
rect 16664 14628 16698 14662
rect 16732 14628 16766 14662
rect 16800 14628 16834 14662
rect 16868 14628 16902 14662
rect 16936 14628 16970 14662
rect 17004 14628 17038 14662
rect 17072 14628 17106 14662
rect 17140 14628 17174 14662
rect 17208 14628 17242 14662
rect 17276 14628 17310 14662
rect 17344 14628 17378 14662
rect 17412 14628 17446 14662
rect 17480 14628 17514 14662
rect 17548 14628 17582 14662
rect 17616 14628 17650 14662
rect 17684 14628 17718 14662
rect 17752 14628 17786 14662
rect 17820 14628 17854 14662
rect 17888 14628 17922 14662
rect 17956 14628 17990 14662
rect 18024 14628 18058 14662
rect 18092 14628 18126 14662
rect 18160 14628 18194 14662
rect 18228 14628 18262 14662
rect 18296 14628 18330 14662
rect 18364 14628 18388 14662
rect 13342 14570 13376 14604
rect 13342 14502 13376 14536
rect 13342 14434 13376 14468
rect 13342 14366 13376 14400
rect 13342 14298 13376 14332
rect 13342 14230 13376 14264
rect 13342 14162 13376 14196
rect 13342 14094 13376 14128
rect 13342 14026 13376 14060
rect 13342 13958 13376 13992
rect 13342 13890 13376 13924
rect 13342 13822 13376 13856
rect 13342 13754 13376 13788
rect 13342 13686 13376 13720
rect 13342 13618 13376 13652
rect 13342 13550 13376 13584
rect 13342 13482 13376 13516
rect 13342 13414 13376 13448
rect 13342 13346 13376 13380
rect 13342 13278 13376 13312
rect 13342 13210 13376 13244
rect 18354 14594 18388 14628
rect 18354 14526 18388 14560
rect 18354 14458 18388 14492
rect 18354 14390 18388 14424
rect 18354 14322 18388 14356
rect 18354 14254 18388 14288
rect 18354 14186 18388 14220
rect 18354 14118 18388 14152
rect 18354 14050 18388 14084
rect 18354 13982 18388 14016
rect 18354 13914 18388 13948
rect 18354 13846 18388 13880
rect 18354 13778 18388 13812
rect 18354 13710 18388 13744
rect 18354 13642 18388 13676
rect 18354 13574 18388 13608
rect 18354 13506 18388 13540
rect 18354 13438 18388 13472
rect 18354 13370 18388 13404
rect 18354 13302 18388 13336
rect 18354 13234 18388 13268
rect 13342 13176 13366 13210
rect 13400 13176 13434 13210
rect 13468 13176 13502 13210
rect 13536 13176 13570 13210
rect 13604 13176 13638 13210
rect 13672 13176 13706 13210
rect 13740 13176 13774 13210
rect 13808 13176 13842 13210
rect 13876 13176 13910 13210
rect 13944 13176 13978 13210
rect 14012 13176 14046 13210
rect 14080 13176 14114 13210
rect 14148 13176 14182 13210
rect 14216 13176 14250 13210
rect 14284 13176 14318 13210
rect 14352 13176 14386 13210
rect 14420 13176 14454 13210
rect 14488 13176 14522 13210
rect 14556 13176 14590 13210
rect 14624 13176 14658 13210
rect 14692 13176 14726 13210
rect 14760 13176 14794 13210
rect 14828 13176 14862 13210
rect 14896 13176 14930 13210
rect 14964 13176 14998 13210
rect 15032 13176 15066 13210
rect 15100 13176 15134 13210
rect 15168 13176 15202 13210
rect 15236 13176 15270 13210
rect 15304 13176 15338 13210
rect 15372 13176 15406 13210
rect 15440 13176 15474 13210
rect 15508 13176 15542 13210
rect 15576 13176 15610 13210
rect 15644 13176 15678 13210
rect 15712 13176 15746 13210
rect 15780 13176 15889 13210
rect 15923 13176 15957 13210
rect 15991 13176 16025 13210
rect 16059 13176 16093 13210
rect 16127 13176 16161 13210
rect 16195 13176 16229 13210
rect 16263 13176 16297 13210
rect 16331 13176 16365 13210
rect 16399 13176 16433 13210
rect 16467 13176 16501 13210
rect 16535 13176 16569 13210
rect 16603 13176 16637 13210
rect 16671 13176 16705 13210
rect 16739 13176 16773 13210
rect 16807 13176 16841 13210
rect 16875 13176 16909 13210
rect 16943 13176 16977 13210
rect 17011 13176 17045 13210
rect 17079 13176 17113 13210
rect 17147 13176 17181 13210
rect 17215 13176 17249 13210
rect 17283 13176 17317 13210
rect 17351 13176 17385 13210
rect 17419 13176 17453 13210
rect 17487 13176 17521 13210
rect 17555 13176 17589 13210
rect 17623 13176 17657 13210
rect 17691 13176 17725 13210
rect 17759 13176 17793 13210
rect 17827 13176 17861 13210
rect 17895 13176 17929 13210
rect 17963 13176 17997 13210
rect 18031 13176 18065 13210
rect 18099 13176 18133 13210
rect 18167 13176 18201 13210
rect 18235 13176 18269 13210
rect 18303 13200 18354 13210
rect 18303 13176 18388 13200
rect 13254 13142 13288 13176
rect 13254 13074 13288 13108
rect 13254 13006 13288 13040
rect 13254 12938 13288 12972
rect 13254 12870 13288 12904
rect 13254 12802 13288 12836
rect 13254 12734 13288 12768
rect 13254 12666 13288 12700
rect 13254 12598 13288 12632
rect 13254 12530 13288 12564
rect 13254 12462 13288 12496
rect 13254 12394 13288 12428
rect 13254 12326 13288 12360
rect 13254 12258 13288 12292
rect 13254 12190 13288 12224
rect 13254 12122 13288 12156
rect 13254 12054 13288 12088
rect 13254 11986 13288 12020
rect 13254 11918 13288 11952
rect 13254 11850 13288 11884
rect 13254 11782 13288 11816
rect 13254 11714 13288 11748
rect 13254 11646 13288 11680
rect 13254 11578 13288 11612
rect 13254 11510 13288 11544
rect 13254 11442 13288 11476
rect 13254 11374 13288 11408
rect 13254 11306 13288 11340
rect 13254 11238 13288 11272
rect 13254 11170 13288 11204
rect 13254 11094 13288 11136
rect 11480 11084 11530 11094
rect 11446 11060 11530 11084
rect 11564 11060 11598 11094
rect 11632 11060 11666 11094
rect 11700 11060 11734 11094
rect 11768 11060 11802 11094
rect 11836 11060 11870 11094
rect 11904 11060 11938 11094
rect 11972 11060 12006 11094
rect 12040 11060 12074 11094
rect 12108 11060 12142 11094
rect 12176 11060 12210 11094
rect 12244 11060 12278 11094
rect 12312 11060 12346 11094
rect 12380 11060 12414 11094
rect 12448 11060 12482 11094
rect 12516 11060 12550 11094
rect 12584 11060 12618 11094
rect 12652 11060 12686 11094
rect 12720 11060 12754 11094
rect 12788 11060 12822 11094
rect 12856 11060 12890 11094
rect 12924 11060 12958 11094
rect 12992 11060 13026 11094
rect 13060 11060 13094 11094
rect 13128 11060 13162 11094
rect 13196 11060 13230 11094
rect 13264 11060 13288 11094
<< nsubdiff >>
rect 9445 37602 9469 37636
rect 9503 37602 9537 37636
rect 9571 37602 9605 37636
rect 9639 37602 9673 37636
rect 9707 37602 9741 37636
rect 9775 37602 9809 37636
rect 9843 37602 9877 37636
rect 9911 37602 9945 37636
rect 9979 37602 10013 37636
rect 10047 37602 10081 37636
rect 10115 37602 10149 37636
rect 10183 37602 10217 37636
rect 10251 37602 10285 37636
rect 10319 37602 10353 37636
rect 10387 37602 10421 37636
rect 10455 37602 10489 37636
rect 10523 37602 10557 37636
rect 10591 37602 10625 37636
rect 10659 37602 10693 37636
rect 10727 37602 10761 37636
rect 10795 37602 10829 37636
rect 10863 37602 10897 37636
rect 10931 37602 10965 37636
rect 10999 37602 11033 37636
rect 11067 37602 11101 37636
rect 11135 37602 11169 37636
rect 11203 37602 11237 37636
rect 11271 37602 11305 37636
rect 11339 37602 11373 37636
rect 11407 37602 11441 37636
rect 11475 37602 11509 37636
rect 11543 37602 11577 37636
rect 11611 37602 11645 37636
rect 11679 37602 11713 37636
rect 11747 37602 11781 37636
rect 11815 37602 11849 37636
rect 11883 37602 11917 37636
rect 11951 37602 11985 37636
rect 12019 37602 12053 37636
rect 12087 37602 12121 37636
rect 12155 37602 12189 37636
rect 12223 37602 12257 37636
rect 12291 37602 12348 37636
rect 12382 37602 12416 37636
rect 12450 37602 12484 37636
rect 12518 37602 12552 37636
rect 12586 37602 12620 37636
rect 12654 37602 12688 37636
rect 12722 37602 12756 37636
rect 12790 37602 12824 37636
rect 12858 37602 12892 37636
rect 12926 37602 12960 37636
rect 12994 37602 13028 37636
rect 13062 37602 13096 37636
rect 13130 37602 13164 37636
rect 13198 37602 13232 37636
rect 13266 37602 13300 37636
rect 13334 37602 13368 37636
rect 13402 37602 13436 37636
rect 13470 37602 13504 37636
rect 13538 37602 13572 37636
rect 13606 37602 13640 37636
rect 13674 37602 13708 37636
rect 13742 37602 13776 37636
rect 13810 37602 13844 37636
rect 13878 37602 13912 37636
rect 13946 37602 13980 37636
rect 14014 37602 14048 37636
rect 14082 37602 14116 37636
rect 14150 37602 14184 37636
rect 14218 37602 14252 37636
rect 14286 37602 14320 37636
rect 14354 37602 14388 37636
rect 14422 37602 14456 37636
rect 14490 37602 14524 37636
rect 14558 37602 14592 37636
rect 14626 37602 14660 37636
rect 14694 37602 14728 37636
rect 14762 37602 14796 37636
rect 14830 37602 14864 37636
rect 14898 37602 14932 37636
rect 14966 37602 15000 37636
rect 15034 37602 15068 37636
rect 15102 37612 15203 37636
rect 15102 37602 15169 37612
rect 9445 37542 9479 37602
rect 15169 37544 15203 37578
rect 9445 37474 9479 37508
rect 9569 37500 10275 37512
rect 9569 37466 9599 37500
rect 9633 37466 9667 37500
rect 9701 37466 9735 37500
rect 9769 37466 9803 37500
rect 9837 37466 9871 37500
rect 9905 37466 9939 37500
rect 9973 37466 10007 37500
rect 10041 37466 10075 37500
rect 10109 37466 10143 37500
rect 10177 37466 10211 37500
rect 10245 37466 10275 37500
rect 9569 37454 10275 37466
rect 10331 37500 14317 37512
rect 10331 37466 10374 37500
rect 10408 37466 10442 37500
rect 10476 37466 10510 37500
rect 10544 37466 10578 37500
rect 10612 37466 10646 37500
rect 10680 37466 10714 37500
rect 10748 37466 10782 37500
rect 10816 37466 10850 37500
rect 10884 37466 10918 37500
rect 10952 37466 11034 37500
rect 11068 37466 11102 37500
rect 11136 37466 11170 37500
rect 11204 37466 11238 37500
rect 11272 37466 11306 37500
rect 11340 37466 11374 37500
rect 11408 37466 11442 37500
rect 11476 37466 11510 37500
rect 11544 37466 11578 37500
rect 11612 37466 11690 37500
rect 11724 37466 11758 37500
rect 11792 37466 11826 37500
rect 11860 37466 11894 37500
rect 11928 37466 11962 37500
rect 11996 37466 12030 37500
rect 12064 37466 12098 37500
rect 12132 37466 12166 37500
rect 12200 37466 12234 37500
rect 12268 37466 12363 37500
rect 12397 37466 12431 37500
rect 12465 37466 12499 37500
rect 12533 37466 12567 37500
rect 12601 37466 12635 37500
rect 12669 37466 12703 37500
rect 12737 37466 12771 37500
rect 12805 37466 12839 37500
rect 12873 37466 12907 37500
rect 12941 37466 13036 37500
rect 13070 37466 13104 37500
rect 13138 37466 13172 37500
rect 13206 37466 13240 37500
rect 13274 37466 13308 37500
rect 13342 37466 13376 37500
rect 13410 37466 13444 37500
rect 13478 37466 13512 37500
rect 13546 37466 13580 37500
rect 13614 37466 13696 37500
rect 13730 37466 13764 37500
rect 13798 37466 13832 37500
rect 13866 37466 13900 37500
rect 13934 37466 13968 37500
rect 14002 37466 14036 37500
rect 14070 37466 14104 37500
rect 14138 37466 14172 37500
rect 14206 37466 14240 37500
rect 14274 37466 14317 37500
rect 10331 37454 14317 37466
rect 15169 37476 15203 37510
rect 9445 37406 9479 37440
rect 15169 37408 15203 37442
rect 9445 37338 9479 37372
rect 9445 37270 9479 37304
rect 9445 37202 9479 37236
rect 9445 37134 9479 37168
rect 9445 37066 9479 37100
rect 9445 36998 9479 37032
rect 9445 36930 9479 36964
rect 9445 36862 9479 36896
rect 9445 36794 9479 36828
rect 9445 36726 9479 36760
rect 9445 36658 9479 36692
rect 9445 36590 9479 36624
rect 9445 36522 9479 36556
rect 9445 36454 9479 36488
rect 9445 36386 9479 36420
rect 9445 36318 9479 36352
rect 9445 36250 9479 36284
rect 9445 36182 9479 36216
rect 9445 36114 9479 36148
rect 9445 36046 9479 36080
rect 15169 37340 15203 37374
rect 15169 37272 15203 37306
rect 15169 37204 15203 37238
rect 15169 37136 15203 37170
rect 15169 37068 15203 37102
rect 15169 37000 15203 37034
rect 15169 36932 15203 36966
rect 15169 36864 15203 36898
rect 15169 36796 15203 36830
rect 15169 36728 15203 36762
rect 15169 36660 15203 36694
rect 15169 36592 15203 36626
rect 15169 36524 15203 36558
rect 15169 36456 15203 36490
rect 15169 36388 15203 36422
rect 15169 36320 15203 36354
rect 15169 36252 15203 36286
rect 15169 36184 15203 36218
rect 15169 36116 15203 36150
rect 15169 36048 15203 36082
rect 9445 35978 9479 36012
rect 15169 35980 15203 36014
rect 9445 35910 9479 35944
rect 9445 35842 9479 35876
rect 9445 35774 9479 35808
rect 9445 35706 9479 35740
rect 9445 35638 9479 35672
rect 9445 35570 9479 35604
rect 9445 35502 9479 35536
rect 9445 35434 9479 35468
rect 9445 35366 9479 35400
rect 9445 35298 9479 35332
rect 9445 35230 9479 35264
rect 9445 35162 9479 35196
rect 9445 35094 9479 35128
rect 9445 35026 9479 35060
rect 9445 34958 9479 34992
rect 9445 34890 9479 34924
rect 9445 34822 9479 34856
rect 9445 34754 9479 34788
rect 6952 34688 6976 34722
rect 7010 34688 7044 34722
rect 7078 34688 7112 34722
rect 7146 34688 7180 34722
rect 7214 34688 7248 34722
rect 7282 34688 7316 34722
rect 7350 34688 7384 34722
rect 7418 34688 7452 34722
rect 7486 34688 7520 34722
rect 7554 34688 7588 34722
rect 7622 34688 7656 34722
rect 7690 34688 7724 34722
rect 7758 34688 7792 34722
rect 7826 34698 7926 34722
rect 7826 34688 7892 34698
rect 6952 34642 6986 34688
rect 6952 34574 6986 34608
rect 6952 34506 6986 34540
rect 6952 34438 6986 34472
rect 6952 34370 6986 34404
rect 6952 34302 6986 34336
rect 6952 34234 6986 34268
rect 6952 34166 6986 34200
rect 6952 34098 6986 34132
rect 6952 34030 6986 34064
rect 6952 33891 6986 33996
rect 6952 33823 6986 33857
rect 6952 33755 6986 33789
rect 6952 33687 6986 33721
rect 6952 33619 6986 33653
rect 6952 33551 6986 33585
rect 6952 33483 6986 33517
rect 6952 33415 6986 33449
rect 6952 33347 6986 33381
rect 6952 33279 6986 33313
rect 7892 34630 7926 34664
rect 7892 34562 7926 34596
rect 7892 34494 7926 34528
rect 7892 34426 7926 34460
rect 9445 34686 9479 34720
rect 9445 34618 9479 34652
rect 15169 35912 15203 35946
rect 15169 35844 15203 35878
rect 15169 35776 15203 35810
rect 15169 35708 15203 35742
rect 15169 35640 15203 35674
rect 15169 35572 15203 35606
rect 15169 35504 15203 35538
rect 15169 35436 15203 35470
rect 15169 35368 15203 35402
rect 15169 35300 15203 35334
rect 15169 35232 15203 35266
rect 15169 35164 15203 35198
rect 15169 35096 15203 35130
rect 15169 35028 15203 35062
rect 15169 34960 15203 34994
rect 15169 34892 15203 34926
rect 15169 34824 15203 34858
rect 15169 34756 15203 34790
rect 15169 34688 15203 34722
rect 15169 34620 15203 34654
rect 9445 34550 9479 34584
rect 15169 34552 15203 34586
rect 9445 34482 9479 34516
rect 15169 34458 15203 34518
rect 9479 34448 9569 34458
rect 9445 34424 9569 34448
rect 9603 34424 9637 34458
rect 9671 34424 9705 34458
rect 9739 34424 9773 34458
rect 9807 34424 9841 34458
rect 9875 34424 9909 34458
rect 9943 34424 9977 34458
rect 10011 34424 10045 34458
rect 10079 34424 10113 34458
rect 10147 34424 10181 34458
rect 10215 34424 10249 34458
rect 10283 34424 10317 34458
rect 10351 34424 10385 34458
rect 10419 34424 10453 34458
rect 10487 34424 10521 34458
rect 10555 34424 10589 34458
rect 10623 34424 10657 34458
rect 10691 34424 10725 34458
rect 10759 34424 10793 34458
rect 10827 34424 10861 34458
rect 10895 34424 10929 34458
rect 10963 34424 10997 34458
rect 11031 34424 11065 34458
rect 11099 34424 11133 34458
rect 11167 34424 11201 34458
rect 11235 34424 11269 34458
rect 11303 34424 11337 34458
rect 11371 34424 11405 34458
rect 11439 34424 11473 34458
rect 11507 34424 11541 34458
rect 11575 34424 11609 34458
rect 11643 34424 11677 34458
rect 11711 34424 11745 34458
rect 11779 34424 11813 34458
rect 11847 34424 11881 34458
rect 11915 34424 11949 34458
rect 11983 34424 12017 34458
rect 12051 34424 12085 34458
rect 12119 34424 12153 34458
rect 12187 34424 12221 34458
rect 12255 34424 12289 34458
rect 12323 34424 12357 34458
rect 12391 34424 12425 34458
rect 12459 34424 12493 34458
rect 12527 34424 12561 34458
rect 12595 34424 12629 34458
rect 12663 34424 12697 34458
rect 12731 34424 12765 34458
rect 12799 34424 12833 34458
rect 12867 34424 12901 34458
rect 12935 34424 12969 34458
rect 13003 34424 13037 34458
rect 13071 34424 13105 34458
rect 13139 34424 13173 34458
rect 13207 34424 13241 34458
rect 13275 34424 13309 34458
rect 13343 34424 13377 34458
rect 13411 34424 13445 34458
rect 13479 34424 13513 34458
rect 13547 34424 13581 34458
rect 13615 34424 13649 34458
rect 13683 34424 13717 34458
rect 13751 34424 13785 34458
rect 13819 34424 13853 34458
rect 13887 34424 13921 34458
rect 13955 34424 13989 34458
rect 14023 34424 14057 34458
rect 14091 34424 14125 34458
rect 14159 34424 14193 34458
rect 14227 34424 14261 34458
rect 14295 34424 14329 34458
rect 14363 34424 14397 34458
rect 14431 34424 14465 34458
rect 14499 34424 14533 34458
rect 14567 34424 14601 34458
rect 14635 34424 14669 34458
rect 14703 34424 14737 34458
rect 14771 34424 14805 34458
rect 14839 34424 14873 34458
rect 14907 34424 14941 34458
rect 14975 34424 15009 34458
rect 15043 34424 15077 34458
rect 15111 34424 15145 34458
rect 15179 34424 15203 34458
rect 15275 37612 15371 37636
rect 15309 37602 15371 37612
rect 15405 37602 15439 37636
rect 15473 37602 15507 37636
rect 15541 37602 15575 37636
rect 15609 37602 15643 37636
rect 15677 37602 15711 37636
rect 15745 37602 15779 37636
rect 15813 37602 15847 37636
rect 15881 37602 15915 37636
rect 15949 37602 15983 37636
rect 16017 37602 16051 37636
rect 16085 37602 16119 37636
rect 16153 37602 16187 37636
rect 16221 37602 16255 37636
rect 16289 37602 16323 37636
rect 16357 37602 16391 37636
rect 16425 37602 16459 37636
rect 16493 37602 16527 37636
rect 16561 37602 16595 37636
rect 16629 37602 16663 37636
rect 16697 37602 16731 37636
rect 16765 37602 16799 37636
rect 16833 37602 16867 37636
rect 16901 37602 16935 37636
rect 16969 37602 17003 37636
rect 17037 37602 17071 37636
rect 17105 37602 17139 37636
rect 17173 37602 17207 37636
rect 17241 37602 17275 37636
rect 17309 37602 17343 37636
rect 17377 37602 17411 37636
rect 17445 37602 17479 37636
rect 17513 37602 17547 37636
rect 17581 37602 17615 37636
rect 17649 37602 17683 37636
rect 17717 37602 17751 37636
rect 17785 37602 17819 37636
rect 17853 37602 17887 37636
rect 17921 37602 17955 37636
rect 17989 37602 18023 37636
rect 18057 37602 18091 37636
rect 18125 37602 18159 37636
rect 18193 37602 18217 37636
rect 15275 37544 15309 37578
rect 15275 37476 15309 37510
rect 15275 37408 15309 37442
rect 15275 37340 15309 37374
rect 15275 37272 15309 37306
rect 15275 37204 15309 37238
rect 15275 37136 15309 37170
rect 15275 37068 15309 37102
rect 15275 37000 15309 37034
rect 15275 36932 15309 36966
rect 15275 36864 15309 36898
rect 15275 36796 15309 36830
rect 15275 36728 15309 36762
rect 15275 36660 15309 36694
rect 15275 36592 15309 36626
rect 15275 36524 15309 36558
rect 15275 36456 15309 36490
rect 15275 36388 15309 36422
rect 15275 36320 15309 36354
rect 15275 36252 15309 36286
rect 15275 36184 15309 36218
rect 15275 36116 15309 36150
rect 15275 36048 15309 36082
rect 15275 35980 15309 36014
rect 15275 35912 15309 35946
rect 15275 35844 15309 35878
rect 15275 35776 15309 35810
rect 15275 35708 15309 35742
rect 15275 35640 15309 35674
rect 15275 35572 15309 35606
rect 15275 35504 15309 35538
rect 15275 35436 15309 35470
rect 15275 35368 15309 35402
rect 15275 35300 15309 35334
rect 15275 35232 15309 35266
rect 15275 35164 15309 35198
rect 15275 35096 15309 35130
rect 15275 35028 15309 35062
rect 15275 34960 15309 34994
rect 15275 34892 15309 34926
rect 15275 34824 15309 34858
rect 15275 34756 15309 34790
rect 15275 34688 15309 34722
rect 15275 34620 15309 34654
rect 15275 34552 15309 34586
rect 15275 34458 15309 34518
rect 18183 37516 18217 37602
rect 18183 37448 18217 37482
rect 18183 37380 18217 37414
rect 18183 37312 18217 37346
rect 18183 37244 18217 37278
rect 18183 37176 18217 37210
rect 18183 37108 18217 37142
rect 18183 37040 18217 37074
rect 18183 36972 18217 37006
rect 18183 36904 18217 36938
rect 18183 36836 18217 36870
rect 18183 36768 18217 36802
rect 18183 36700 18217 36734
rect 18183 36632 18217 36666
rect 18183 36564 18217 36598
rect 18183 36496 18217 36530
rect 18183 36428 18217 36462
rect 18183 36360 18217 36394
rect 18183 36292 18217 36326
rect 18183 36224 18217 36258
rect 18183 36156 18217 36190
rect 18183 36088 18217 36122
rect 18183 35978 18217 36054
rect 18183 35910 18217 35944
rect 18183 35842 18217 35876
rect 18183 35774 18217 35808
rect 18183 35706 18217 35740
rect 18183 35638 18217 35672
rect 18183 35570 18217 35604
rect 18183 35502 18217 35536
rect 18183 35434 18217 35468
rect 18183 35366 18217 35400
rect 18183 35298 18217 35332
rect 18183 35230 18217 35264
rect 18183 35162 18217 35196
rect 18183 35094 18217 35128
rect 18183 35026 18217 35060
rect 18183 34958 18217 34992
rect 18183 34890 18217 34924
rect 18183 34822 18217 34856
rect 18183 34754 18217 34788
rect 18183 34686 18217 34720
rect 18183 34618 18217 34652
rect 18183 34550 18217 34584
rect 18183 34482 18217 34516
rect 15275 34424 15299 34458
rect 15333 34424 15367 34458
rect 15401 34424 15435 34458
rect 15469 34424 15503 34458
rect 15537 34424 15571 34458
rect 15605 34424 15639 34458
rect 15673 34424 15707 34458
rect 15741 34424 15775 34458
rect 15809 34424 15843 34458
rect 15877 34424 15911 34458
rect 15945 34424 15979 34458
rect 16013 34424 16047 34458
rect 16081 34424 16115 34458
rect 16149 34424 16183 34458
rect 16217 34424 16251 34458
rect 16285 34424 16319 34458
rect 16353 34424 16387 34458
rect 16421 34424 16455 34458
rect 16489 34424 16523 34458
rect 16557 34424 16591 34458
rect 16625 34424 16659 34458
rect 16693 34424 16727 34458
rect 16761 34424 16795 34458
rect 16829 34424 16863 34458
rect 16897 34424 16931 34458
rect 16965 34424 16999 34458
rect 17033 34424 17067 34458
rect 17101 34424 17135 34458
rect 17169 34424 17203 34458
rect 17237 34424 17271 34458
rect 17305 34424 17339 34458
rect 17373 34424 17407 34458
rect 17441 34424 17475 34458
rect 17509 34424 17543 34458
rect 17577 34424 17611 34458
rect 17645 34424 17679 34458
rect 17713 34424 17747 34458
rect 17781 34424 17815 34458
rect 17849 34424 17883 34458
rect 17917 34424 17951 34458
rect 17985 34424 18019 34458
rect 18053 34424 18087 34458
rect 18121 34448 18183 34458
rect 18121 34424 18217 34448
rect 18289 37612 18362 37636
rect 18323 37602 18362 37612
rect 18396 37602 18430 37636
rect 18464 37602 18498 37636
rect 18532 37602 18566 37636
rect 18600 37602 18634 37636
rect 18668 37602 18702 37636
rect 18736 37602 18770 37636
rect 18804 37602 18838 37636
rect 18872 37602 18906 37636
rect 18940 37602 18974 37636
rect 19008 37602 19042 37636
rect 19076 37602 19110 37636
rect 19144 37602 19178 37636
rect 19212 37602 19246 37636
rect 19280 37602 19314 37636
rect 19348 37602 19382 37636
rect 19416 37602 19450 37636
rect 19484 37602 19518 37636
rect 19552 37602 19586 37636
rect 19620 37602 19654 37636
rect 19688 37602 19722 37636
rect 19756 37602 19790 37636
rect 19824 37602 19858 37636
rect 19892 37602 19926 37636
rect 19960 37602 19994 37636
rect 20028 37602 20062 37636
rect 20096 37602 20130 37636
rect 20164 37602 20198 37636
rect 20232 37602 20266 37636
rect 20300 37602 20334 37636
rect 20368 37602 20402 37636
rect 20436 37602 20470 37636
rect 20504 37602 20538 37636
rect 20572 37602 20606 37636
rect 20640 37602 20674 37636
rect 20708 37602 20742 37636
rect 20776 37602 20810 37636
rect 20844 37602 20878 37636
rect 20912 37602 20946 37636
rect 20980 37602 21014 37636
rect 21048 37602 21145 37636
rect 21179 37602 21213 37636
rect 21247 37602 21281 37636
rect 21315 37602 21349 37636
rect 21383 37602 21417 37636
rect 21451 37602 21485 37636
rect 21519 37602 21553 37636
rect 21587 37602 21621 37636
rect 21655 37602 21689 37636
rect 21723 37602 21757 37636
rect 21791 37602 21825 37636
rect 21859 37602 21893 37636
rect 21927 37602 21961 37636
rect 21995 37602 22029 37636
rect 22063 37602 22097 37636
rect 22131 37602 22165 37636
rect 22199 37602 22233 37636
rect 22267 37602 22301 37636
rect 22335 37602 22369 37636
rect 22403 37602 22437 37636
rect 22471 37602 22505 37636
rect 22539 37602 22573 37636
rect 22607 37602 22641 37636
rect 22675 37602 22709 37636
rect 22743 37602 22777 37636
rect 22811 37602 22845 37636
rect 22879 37602 22913 37636
rect 22947 37602 22981 37636
rect 23015 37602 23049 37636
rect 23083 37602 23117 37636
rect 23151 37602 23185 37636
rect 23219 37602 23253 37636
rect 23287 37602 23321 37636
rect 23355 37602 23389 37636
rect 23423 37602 23457 37636
rect 23491 37602 23525 37636
rect 23559 37602 23593 37636
rect 23627 37602 23661 37636
rect 23695 37602 23729 37636
rect 23763 37602 23797 37636
rect 23831 37602 23855 37636
rect 18289 37544 18323 37578
rect 18289 37476 18323 37510
rect 23821 37542 23855 37602
rect 18289 37408 18323 37442
rect 19087 37482 23057 37494
rect 19087 37448 19143 37482
rect 19177 37448 19211 37482
rect 19245 37448 19279 37482
rect 19313 37448 19347 37482
rect 19381 37448 19415 37482
rect 19449 37448 19483 37482
rect 19517 37448 19551 37482
rect 19585 37448 19619 37482
rect 19653 37448 19687 37482
rect 19721 37448 19816 37482
rect 19850 37448 19884 37482
rect 19918 37448 19952 37482
rect 19986 37448 20020 37482
rect 20054 37448 20088 37482
rect 20122 37448 20156 37482
rect 20190 37448 20224 37482
rect 20258 37448 20292 37482
rect 20326 37448 20360 37482
rect 20394 37448 20489 37482
rect 20523 37448 20557 37482
rect 20591 37448 20625 37482
rect 20659 37448 20693 37482
rect 20727 37448 20761 37482
rect 20795 37448 20829 37482
rect 20863 37448 20897 37482
rect 20931 37448 20965 37482
rect 20999 37448 21094 37482
rect 21128 37448 21162 37482
rect 21196 37448 21230 37482
rect 21264 37448 21298 37482
rect 21332 37448 21366 37482
rect 21400 37448 21434 37482
rect 21468 37448 21502 37482
rect 21536 37448 21570 37482
rect 21604 37448 21638 37482
rect 21672 37448 21767 37482
rect 21801 37448 21835 37482
rect 21869 37448 21903 37482
rect 21937 37448 21971 37482
rect 22005 37448 22039 37482
rect 22073 37448 22107 37482
rect 22141 37448 22175 37482
rect 22209 37448 22243 37482
rect 22277 37448 22311 37482
rect 22345 37448 22440 37482
rect 22474 37448 22508 37482
rect 22542 37448 22576 37482
rect 22610 37448 22644 37482
rect 22678 37448 22712 37482
rect 22746 37448 22780 37482
rect 22814 37448 22848 37482
rect 22882 37448 22916 37482
rect 22950 37448 22984 37482
rect 23018 37448 23057 37482
rect 19087 37436 23057 37448
rect 23821 37474 23855 37508
rect 23821 37406 23855 37440
rect 18289 37340 18323 37374
rect 18289 37272 18323 37306
rect 18289 37204 18323 37238
rect 18289 37136 18323 37170
rect 18289 37068 18323 37102
rect 18289 37000 18323 37034
rect 18289 36932 18323 36966
rect 18289 36864 18323 36898
rect 18289 36796 18323 36830
rect 18289 36728 18323 36762
rect 18289 36660 18323 36694
rect 18289 36592 18323 36626
rect 18289 36524 18323 36558
rect 18289 36456 18323 36490
rect 18289 36388 18323 36422
rect 18289 36320 18323 36354
rect 18289 36252 18323 36286
rect 18289 36184 18323 36218
rect 18289 36116 18323 36150
rect 18289 36048 18323 36082
rect 23821 37338 23855 37372
rect 23821 37270 23855 37304
rect 23821 37202 23855 37236
rect 23821 37134 23855 37168
rect 23821 37066 23855 37100
rect 23821 36998 23855 37032
rect 23821 36930 23855 36964
rect 23821 36862 23855 36896
rect 23821 36794 23855 36828
rect 23821 36726 23855 36760
rect 23821 36658 23855 36692
rect 23821 36590 23855 36624
rect 23821 36522 23855 36556
rect 23821 36454 23855 36488
rect 23821 36386 23855 36420
rect 23821 36318 23855 36352
rect 23821 36250 23855 36284
rect 23821 36182 23855 36216
rect 23821 36114 23855 36148
rect 23821 36046 23855 36080
rect 18289 35980 18323 36014
rect 18289 35912 18323 35946
rect 18289 35844 18323 35878
rect 18289 35776 18323 35810
rect 18289 35708 18323 35742
rect 18289 35640 18323 35674
rect 18289 35572 18323 35606
rect 18289 35504 18323 35538
rect 18289 35436 18323 35470
rect 18289 35368 18323 35402
rect 18289 35300 18323 35334
rect 18289 35232 18323 35266
rect 18289 35164 18323 35198
rect 18289 35096 18323 35130
rect 18289 35028 18323 35062
rect 18289 34960 18323 34994
rect 18289 34892 18323 34926
rect 18289 34824 18323 34858
rect 18289 34756 18323 34790
rect 18289 34688 18323 34722
rect 18289 34620 18323 34654
rect 18289 34552 18323 34586
rect 18289 34458 18323 34518
rect 23821 35978 23855 36012
rect 23821 35910 23855 35944
rect 23821 35842 23855 35876
rect 23821 35774 23855 35808
rect 23821 35706 23855 35740
rect 23821 35638 23855 35672
rect 23821 35570 23855 35604
rect 23821 35502 23855 35536
rect 23821 35434 23855 35468
rect 23821 35366 23855 35400
rect 23821 35298 23855 35332
rect 23821 35230 23855 35264
rect 23821 35162 23855 35196
rect 23821 35094 23855 35128
rect 23821 35026 23855 35060
rect 23821 34958 23855 34992
rect 23821 34890 23855 34924
rect 23821 34822 23855 34856
rect 23821 34754 23855 34788
rect 23821 34686 23855 34720
rect 23821 34618 23855 34652
rect 23821 34550 23855 34584
rect 23821 34482 23855 34516
rect 18289 34424 18313 34458
rect 18347 34424 18381 34458
rect 18415 34424 18449 34458
rect 18483 34424 18517 34458
rect 18551 34424 18585 34458
rect 18619 34424 18653 34458
rect 18687 34424 18721 34458
rect 18755 34424 18789 34458
rect 18823 34424 18857 34458
rect 18891 34424 18925 34458
rect 18959 34424 18993 34458
rect 19027 34424 19061 34458
rect 19095 34424 19129 34458
rect 19163 34424 19197 34458
rect 19231 34424 19265 34458
rect 19299 34424 19333 34458
rect 19367 34424 19401 34458
rect 19435 34424 19469 34458
rect 19503 34424 19537 34458
rect 19571 34424 19605 34458
rect 19639 34424 19673 34458
rect 19707 34424 19741 34458
rect 19775 34424 19809 34458
rect 19843 34424 19877 34458
rect 19911 34424 19945 34458
rect 19979 34424 20013 34458
rect 20047 34424 20081 34458
rect 20115 34424 20149 34458
rect 20183 34424 20217 34458
rect 20251 34424 20285 34458
rect 20319 34424 20353 34458
rect 20387 34424 20421 34458
rect 20455 34424 20489 34458
rect 20523 34424 20557 34458
rect 20591 34424 20625 34458
rect 20659 34424 20693 34458
rect 20727 34424 20761 34458
rect 20795 34424 20829 34458
rect 20863 34424 20897 34458
rect 20931 34424 20965 34458
rect 20999 34424 21033 34458
rect 21067 34424 21101 34458
rect 21135 34424 21169 34458
rect 21203 34424 21237 34458
rect 21271 34424 21305 34458
rect 21339 34424 21373 34458
rect 21407 34424 21441 34458
rect 21475 34424 21509 34458
rect 21543 34424 21577 34458
rect 21611 34424 21645 34458
rect 21679 34424 21713 34458
rect 21747 34424 21781 34458
rect 21815 34424 21849 34458
rect 21883 34424 21917 34458
rect 21951 34424 21985 34458
rect 22019 34424 22053 34458
rect 22087 34424 22121 34458
rect 22155 34424 22189 34458
rect 22223 34424 22257 34458
rect 22291 34424 22325 34458
rect 22359 34424 22393 34458
rect 22427 34424 22461 34458
rect 22495 34424 22529 34458
rect 22563 34424 22597 34458
rect 22631 34424 22665 34458
rect 22699 34424 22733 34458
rect 22767 34424 22801 34458
rect 22835 34424 22869 34458
rect 22903 34424 22937 34458
rect 22971 34424 23005 34458
rect 23039 34424 23073 34458
rect 23107 34424 23141 34458
rect 23175 34424 23209 34458
rect 23243 34424 23277 34458
rect 23311 34424 23345 34458
rect 23379 34424 23413 34458
rect 23447 34424 23481 34458
rect 23515 34424 23549 34458
rect 23583 34424 23617 34458
rect 23651 34424 23685 34458
rect 23719 34424 23753 34458
rect 23787 34448 23821 34458
rect 23787 34424 23855 34448
rect 7892 34358 7926 34392
rect 7892 34290 7926 34324
rect 7892 34222 7926 34256
rect 7892 34154 7926 34188
rect 7892 34086 7926 34120
rect 7892 34018 7926 34052
rect 7892 33950 7926 33984
rect 7892 33882 7926 33916
rect 7892 33814 7926 33848
rect 7892 33746 7926 33780
rect 7892 33678 7926 33712
rect 9445 34318 9469 34352
rect 9503 34318 9537 34352
rect 9571 34318 9605 34352
rect 9639 34318 9673 34352
rect 9707 34318 9741 34352
rect 9775 34318 9809 34352
rect 9843 34318 9877 34352
rect 9911 34318 9945 34352
rect 9979 34318 10013 34352
rect 10047 34318 10081 34352
rect 10115 34318 10149 34352
rect 10183 34318 10217 34352
rect 10251 34318 10285 34352
rect 10319 34318 10353 34352
rect 10387 34318 10421 34352
rect 10455 34318 10489 34352
rect 10523 34318 10637 34352
rect 10671 34318 10705 34352
rect 10739 34318 10773 34352
rect 10807 34318 10841 34352
rect 10875 34318 10909 34352
rect 10943 34318 10977 34352
rect 11011 34318 11045 34352
rect 11079 34318 11113 34352
rect 11147 34318 11181 34352
rect 11215 34318 11249 34352
rect 11283 34318 11317 34352
rect 11351 34318 11385 34352
rect 11419 34318 11453 34352
rect 11487 34318 11521 34352
rect 11555 34318 11589 34352
rect 11623 34318 11657 34352
rect 11691 34328 11781 34352
rect 15203 34351 15227 34352
rect 11691 34318 11747 34328
rect 9445 34278 9479 34318
rect 9445 34210 9479 34244
rect 11747 34260 11781 34294
rect 11747 34192 11781 34226
rect 9445 34142 9479 34176
rect 9445 34074 9479 34108
rect 11747 34124 11781 34158
rect 9445 34006 9479 34040
rect 9445 33938 9479 33972
rect 9445 33870 9479 33904
rect 9445 33802 9479 33836
rect 9445 33734 9479 33768
rect 9445 33666 9479 33700
rect 7892 33610 7926 33644
rect 9445 33598 9479 33632
rect 7892 33542 7926 33576
rect 7892 33474 7926 33508
rect 9445 33530 9479 33564
rect 9655 34054 9713 34099
rect 9655 34020 9667 34054
rect 9701 34020 9713 34054
rect 9655 33986 9713 34020
rect 9655 33952 9667 33986
rect 9701 33952 9713 33986
rect 9655 33918 9713 33952
rect 9655 33884 9667 33918
rect 9701 33884 9713 33918
rect 9655 33850 9713 33884
rect 9655 33816 9667 33850
rect 9701 33816 9713 33850
rect 9655 33782 9713 33816
rect 9655 33748 9667 33782
rect 9701 33748 9713 33782
rect 9655 33714 9713 33748
rect 9655 33680 9667 33714
rect 9701 33680 9713 33714
rect 9655 33646 9713 33680
rect 9655 33612 9667 33646
rect 9701 33612 9713 33646
rect 9655 33578 9713 33612
rect 9655 33544 9667 33578
rect 9701 33544 9713 33578
rect 9655 33499 9713 33544
rect 11513 34054 11571 34099
rect 11513 34020 11525 34054
rect 11559 34020 11571 34054
rect 11513 33986 11571 34020
rect 11513 33952 11525 33986
rect 11559 33952 11571 33986
rect 11513 33918 11571 33952
rect 11513 33884 11525 33918
rect 11559 33884 11571 33918
rect 11513 33850 11571 33884
rect 11513 33816 11525 33850
rect 11559 33816 11571 33850
rect 11513 33782 11571 33816
rect 11513 33748 11525 33782
rect 11559 33748 11571 33782
rect 11513 33714 11571 33748
rect 11513 33680 11525 33714
rect 11559 33680 11571 33714
rect 11513 33646 11571 33680
rect 11513 33612 11525 33646
rect 11559 33612 11571 33646
rect 11513 33578 11571 33612
rect 11513 33544 11525 33578
rect 11559 33544 11571 33578
rect 11513 33499 11571 33544
rect 11747 34056 11781 34090
rect 11747 33988 11781 34022
rect 11747 33920 11781 33954
rect 11747 33852 11781 33886
rect 11747 33784 11781 33818
rect 11747 33716 11781 33750
rect 11747 33648 11781 33682
rect 11747 33580 11781 33614
rect 11747 33512 11781 33546
rect 9445 33462 9479 33496
rect 7892 33406 7926 33440
rect 7892 33338 7926 33372
rect 7892 33255 7926 33304
rect 6986 33245 7052 33255
rect 6952 33221 7052 33245
rect 7086 33221 7120 33255
rect 7154 33221 7188 33255
rect 7222 33221 7256 33255
rect 7290 33221 7324 33255
rect 7358 33221 7392 33255
rect 7426 33221 7460 33255
rect 7494 33221 7528 33255
rect 7562 33221 7596 33255
rect 7630 33221 7664 33255
rect 7698 33221 7732 33255
rect 7766 33221 7800 33255
rect 7834 33221 7868 33255
rect 7902 33221 7926 33255
rect 9445 33394 9479 33428
rect 11747 33444 11781 33478
rect 9445 33326 9479 33360
rect 9445 33258 9479 33292
rect 11747 33376 11781 33410
rect 11747 33308 11781 33342
rect 11747 33234 11781 33274
rect 9479 33224 9547 33234
rect 9445 33200 9547 33224
rect 9581 33200 9615 33234
rect 9649 33200 9683 33234
rect 9717 33200 9751 33234
rect 9785 33200 9819 33234
rect 9853 33200 9887 33234
rect 9921 33200 9955 33234
rect 9989 33200 10023 33234
rect 10057 33200 10091 33234
rect 10125 33200 10159 33234
rect 10193 33200 10227 33234
rect 10261 33200 10295 33234
rect 10329 33200 10363 33234
rect 10397 33200 10431 33234
rect 10465 33200 10499 33234
rect 10533 33200 10567 33234
rect 10601 33200 10635 33234
rect 10669 33200 10703 33234
rect 10737 33200 10771 33234
rect 10805 33200 10839 33234
rect 10873 33200 10907 33234
rect 10941 33200 10975 33234
rect 11009 33200 11043 33234
rect 11077 33200 11111 33234
rect 11145 33200 11179 33234
rect 11213 33200 11247 33234
rect 11281 33200 11315 33234
rect 11349 33200 11383 33234
rect 11417 33200 11451 33234
rect 11485 33200 11519 33234
rect 11553 33200 11587 33234
rect 11621 33200 11655 33234
rect 11689 33200 11723 33234
rect 11757 33200 11781 33234
rect 11853 34316 11877 34350
rect 11911 34316 11945 34350
rect 11979 34316 12013 34350
rect 12047 34316 12081 34350
rect 12115 34316 12149 34350
rect 12183 34316 12217 34350
rect 12251 34316 12285 34350
rect 12319 34316 12353 34350
rect 12387 34316 12421 34350
rect 12455 34316 12489 34350
rect 12523 34316 12557 34350
rect 12591 34316 12625 34350
rect 12659 34316 12693 34350
rect 12727 34316 12761 34350
rect 12795 34326 12919 34350
rect 12795 34316 12885 34326
rect 11853 34241 11887 34316
rect 12885 34258 12919 34292
rect 11853 34173 11887 34207
rect 11955 34238 12773 34250
rect 11955 34204 12002 34238
rect 12036 34204 12070 34238
rect 12104 34204 12138 34238
rect 12172 34204 12262 34238
rect 12296 34204 12330 34238
rect 12364 34204 12398 34238
rect 12432 34204 12505 34238
rect 12539 34204 12573 34238
rect 12607 34204 12641 34238
rect 12675 34204 12709 34238
rect 12743 34204 12773 34238
rect 11955 34192 12773 34204
rect 12885 34190 12919 34224
rect 11853 34105 11887 34139
rect 11853 34037 11887 34071
rect 11853 33969 11887 34003
rect 11853 33901 11887 33935
rect 11853 33833 11887 33867
rect 11853 33734 11887 33799
rect 11853 33666 11887 33700
rect 11853 33598 11887 33632
rect 11853 33530 11887 33564
rect 11853 33462 11887 33496
rect 11853 33394 11887 33428
rect 12885 34122 12919 34156
rect 12885 34054 12919 34088
rect 12885 33986 12919 34020
rect 12885 33918 12919 33952
rect 12885 33850 12919 33884
rect 12885 33782 12919 33816
rect 12885 33714 12919 33748
rect 12885 33646 12919 33680
rect 12885 33578 12919 33612
rect 12885 33510 12919 33544
rect 12885 33442 12919 33476
rect 11853 33326 11887 33360
rect 12885 33374 12919 33408
rect 11853 33258 11887 33292
rect 12885 33306 12919 33340
rect 12885 33234 12919 33272
rect 11887 33224 11977 33234
rect 11853 33200 11977 33224
rect 12011 33200 12045 33234
rect 12079 33200 12113 33234
rect 12147 33200 12181 33234
rect 12215 33200 12249 33234
rect 12283 33200 12317 33234
rect 12351 33200 12385 33234
rect 12419 33200 12453 33234
rect 12487 33200 12521 33234
rect 12555 33200 12589 33234
rect 12623 33200 12657 33234
rect 12691 33200 12725 33234
rect 12759 33200 12793 33234
rect 12827 33200 12861 33234
rect 12895 33200 12919 33234
rect 12991 34317 13015 34351
rect 13049 34317 13083 34351
rect 13117 34317 13151 34351
rect 13185 34317 13219 34351
rect 13253 34317 13287 34351
rect 13321 34317 13355 34351
rect 13389 34317 13423 34351
rect 13457 34317 13491 34351
rect 13525 34317 13559 34351
rect 13593 34317 13627 34351
rect 13661 34317 13695 34351
rect 13729 34317 13763 34351
rect 13797 34317 13831 34351
rect 13865 34317 13899 34351
rect 13933 34317 13967 34351
rect 14001 34317 14035 34351
rect 14069 34317 14103 34351
rect 14137 34317 14171 34351
rect 14205 34317 14239 34351
rect 14273 34317 14307 34351
rect 14341 34317 14375 34351
rect 14409 34317 14443 34351
rect 14477 34317 14511 34351
rect 14545 34317 14579 34351
rect 14613 34317 14647 34351
rect 14681 34317 14715 34351
rect 14749 34317 14783 34351
rect 14817 34317 14851 34351
rect 14885 34317 14919 34351
rect 14953 34317 14987 34351
rect 15021 34317 15055 34351
rect 15089 34317 15123 34351
rect 15157 34318 15227 34351
rect 15261 34318 15295 34352
rect 15329 34318 15363 34352
rect 15397 34318 15431 34352
rect 15465 34318 15499 34352
rect 15533 34318 15567 34352
rect 15601 34318 15635 34352
rect 15669 34318 15703 34352
rect 15737 34318 15771 34352
rect 15805 34318 15839 34352
rect 15873 34318 15907 34352
rect 15941 34318 15975 34352
rect 16009 34318 16043 34352
rect 16077 34328 16193 34352
rect 16077 34318 16159 34328
rect 15157 34317 15237 34318
rect 12991 34278 13025 34317
rect 12991 34210 13025 34244
rect 16159 34260 16193 34294
rect 12991 34142 13025 34176
rect 13089 34220 13795 34232
rect 13089 34186 13119 34220
rect 13153 34186 13187 34220
rect 13221 34186 13255 34220
rect 13289 34186 13323 34220
rect 13357 34186 13391 34220
rect 13425 34186 13459 34220
rect 13493 34186 13527 34220
rect 13561 34186 13595 34220
rect 13629 34186 13663 34220
rect 13697 34186 13731 34220
rect 13765 34186 13795 34220
rect 13089 34174 13795 34186
rect 13867 34220 14565 34232
rect 13867 34186 13893 34220
rect 13927 34186 13961 34220
rect 13995 34186 14029 34220
rect 14063 34186 14097 34220
rect 14131 34186 14165 34220
rect 14199 34186 14233 34220
rect 14267 34186 14301 34220
rect 14335 34186 14369 34220
rect 14403 34186 14437 34220
rect 14471 34186 14505 34220
rect 14539 34186 14565 34220
rect 13867 34174 14565 34186
rect 16159 34192 16193 34226
rect 12991 34074 13025 34108
rect 16159 34124 16193 34158
rect 12991 34006 13025 34040
rect 12991 33938 13025 33972
rect 12991 33870 13025 33904
rect 12991 33802 13025 33836
rect 12991 33734 13025 33768
rect 12991 33666 13025 33700
rect 12991 33598 13025 33632
rect 12991 33530 13025 33564
rect 12991 33462 13025 33496
rect 16159 34056 16193 34090
rect 16159 33988 16193 34022
rect 16159 33920 16193 33954
rect 16159 33852 16193 33886
rect 16159 33784 16193 33818
rect 16159 33716 16193 33750
rect 16159 33648 16193 33682
rect 16159 33580 16193 33614
rect 16159 33512 16193 33546
rect 16159 33444 16193 33478
rect 12991 33394 13025 33428
rect 12991 33326 13025 33360
rect 16159 33376 16193 33410
rect 12991 33258 13025 33292
rect 16159 33308 16193 33342
rect 16159 33234 16193 33274
rect 13025 33224 13106 33234
rect 12991 33200 13106 33224
rect 13140 33200 13174 33234
rect 13208 33200 13242 33234
rect 13276 33200 13310 33234
rect 13344 33200 13378 33234
rect 13412 33200 13446 33234
rect 13480 33200 13514 33234
rect 13548 33200 13582 33234
rect 13616 33200 13650 33234
rect 13684 33200 13718 33234
rect 13752 33200 13786 33234
rect 13820 33200 13854 33234
rect 13888 33200 13922 33234
rect 13956 33200 13990 33234
rect 14024 33200 14058 33234
rect 14092 33200 14126 33234
rect 14160 33200 14194 33234
rect 14228 33200 14262 33234
rect 14296 33200 14330 33234
rect 14364 33200 14398 33234
rect 14432 33200 14466 33234
rect 14500 33200 14534 33234
rect 14568 33200 14639 33234
rect 14673 33200 14707 33234
rect 14741 33200 14775 33234
rect 14809 33200 14843 33234
rect 14877 33200 14911 33234
rect 14945 33200 14979 33234
rect 15013 33200 15047 33234
rect 15081 33200 15115 33234
rect 15149 33200 15183 33234
rect 15217 33200 15251 33234
rect 15285 33200 15319 33234
rect 15353 33200 15387 33234
rect 15421 33200 15455 33234
rect 15489 33200 15523 33234
rect 15557 33200 15591 33234
rect 15625 33200 15659 33234
rect 15693 33200 15727 33234
rect 15761 33200 15795 33234
rect 15829 33200 15863 33234
rect 15897 33200 15931 33234
rect 15965 33200 15999 33234
rect 16033 33200 16067 33234
rect 16101 33200 16135 33234
rect 16169 33200 16193 33234
rect 11457 19226 11481 19260
rect 11515 19226 11549 19260
rect 11583 19226 11617 19260
rect 11651 19226 11685 19260
rect 11719 19226 11753 19260
rect 11787 19226 11821 19260
rect 11855 19226 11889 19260
rect 11923 19226 11957 19260
rect 11991 19226 12025 19260
rect 12059 19226 12093 19260
rect 12127 19226 12161 19260
rect 12195 19226 12229 19260
rect 12263 19226 12297 19260
rect 12331 19226 12365 19260
rect 12399 19226 12433 19260
rect 12467 19226 12501 19260
rect 12535 19226 12569 19260
rect 12603 19226 12637 19260
rect 12671 19226 12705 19260
rect 12739 19226 12773 19260
rect 12807 19226 12841 19260
rect 12875 19226 12909 19260
rect 12943 19226 12977 19260
rect 13011 19226 13045 19260
rect 13079 19226 13113 19260
rect 13147 19226 13181 19260
rect 13215 19226 13249 19260
rect 13283 19226 13317 19260
rect 13351 19226 13385 19260
rect 13419 19226 13453 19260
rect 13487 19226 13521 19260
rect 13555 19226 13589 19260
rect 13623 19226 13657 19260
rect 13691 19226 13725 19260
rect 13759 19226 13793 19260
rect 13827 19226 13861 19260
rect 13895 19226 13929 19260
rect 13963 19226 13997 19260
rect 14031 19226 14065 19260
rect 14099 19226 14133 19260
rect 14167 19226 14201 19260
rect 14235 19226 14269 19260
rect 14303 19226 14360 19260
rect 14394 19226 14428 19260
rect 14462 19226 14496 19260
rect 14530 19226 14564 19260
rect 14598 19226 14632 19260
rect 14666 19226 14700 19260
rect 14734 19226 14768 19260
rect 14802 19226 14836 19260
rect 14870 19226 14904 19260
rect 14938 19226 14972 19260
rect 15006 19226 15040 19260
rect 15074 19226 15108 19260
rect 15142 19226 15176 19260
rect 15210 19226 15244 19260
rect 15278 19226 15312 19260
rect 15346 19226 15380 19260
rect 15414 19226 15448 19260
rect 15482 19226 15516 19260
rect 15550 19226 15584 19260
rect 15618 19226 15652 19260
rect 15686 19226 15720 19260
rect 15754 19226 15788 19260
rect 15822 19226 15856 19260
rect 15890 19226 15924 19260
rect 15958 19226 15992 19260
rect 16026 19226 16060 19260
rect 16094 19226 16128 19260
rect 16162 19226 16196 19260
rect 16230 19226 16264 19260
rect 16298 19226 16332 19260
rect 16366 19226 16400 19260
rect 16434 19226 16468 19260
rect 16502 19226 16536 19260
rect 16570 19226 16604 19260
rect 16638 19226 16672 19260
rect 16706 19226 16740 19260
rect 16774 19226 16808 19260
rect 16842 19226 16876 19260
rect 16910 19226 16944 19260
rect 16978 19226 17012 19260
rect 17046 19226 17080 19260
rect 17114 19236 17215 19260
rect 17114 19226 17181 19236
rect 11457 19166 11491 19226
rect 11457 19098 11491 19132
rect 11457 19030 11491 19064
rect 11457 18962 11491 18996
rect 11457 18894 11491 18928
rect 11457 18826 11491 18860
rect 11457 18758 11491 18792
rect 11457 18690 11491 18724
rect 11457 18622 11491 18656
rect 11457 18554 11491 18588
rect 11457 18486 11491 18520
rect 11457 18418 11491 18452
rect 11457 18350 11491 18384
rect 11457 18282 11491 18316
rect 11457 18214 11491 18248
rect 11457 18146 11491 18180
rect 11457 18078 11491 18112
rect 11457 18010 11491 18044
rect 11457 17942 11491 17976
rect 11457 17874 11491 17908
rect 11457 17806 11491 17840
rect 11457 17738 11491 17772
rect 11457 17670 11491 17704
rect 17181 19168 17215 19202
rect 17181 19100 17215 19134
rect 17181 19032 17215 19066
rect 17181 18964 17215 18998
rect 17181 18896 17215 18930
rect 17181 18828 17215 18862
rect 17181 18760 17215 18794
rect 17181 18692 17215 18726
rect 17181 18624 17215 18658
rect 17181 18556 17215 18590
rect 17181 18488 17215 18522
rect 17181 18420 17215 18454
rect 17181 18352 17215 18386
rect 17181 18284 17215 18318
rect 17181 18216 17215 18250
rect 17181 18148 17215 18182
rect 17181 18080 17215 18114
rect 17181 18012 17215 18046
rect 17181 17944 17215 17978
rect 17181 17876 17215 17910
rect 17181 17808 17215 17842
rect 17181 17740 17215 17774
rect 17181 17672 17215 17706
rect 11457 17602 11491 17636
rect 11457 17534 11491 17568
rect 11457 17466 11491 17500
rect 11457 17398 11491 17432
rect 11457 17330 11491 17364
rect 11457 17262 11491 17296
rect 11457 17194 11491 17228
rect 11457 17126 11491 17160
rect 11457 17058 11491 17092
rect 11457 16990 11491 17024
rect 11457 16922 11491 16956
rect 11457 16854 11491 16888
rect 11457 16786 11491 16820
rect 11457 16718 11491 16752
rect 11457 16650 11491 16684
rect 11457 16582 11491 16616
rect 11457 16514 11491 16548
rect 11457 16446 11491 16480
rect 11457 16378 11491 16412
rect 8964 16312 8988 16346
rect 9022 16312 9056 16346
rect 9090 16312 9124 16346
rect 9158 16312 9192 16346
rect 9226 16312 9260 16346
rect 9294 16312 9328 16346
rect 9362 16312 9396 16346
rect 9430 16312 9464 16346
rect 9498 16312 9532 16346
rect 9566 16312 9600 16346
rect 9634 16312 9668 16346
rect 9702 16312 9736 16346
rect 9770 16312 9804 16346
rect 9838 16322 9938 16346
rect 9838 16312 9904 16322
rect 8964 16266 8998 16312
rect 8964 16198 8998 16232
rect 8964 16130 8998 16164
rect 8964 16062 8998 16096
rect 8964 15994 8998 16028
rect 8964 15926 8998 15960
rect 8964 15858 8998 15892
rect 8964 15790 8998 15824
rect 8964 15722 8998 15756
rect 8964 15654 8998 15688
rect 8964 15515 8998 15620
rect 8964 15447 8998 15481
rect 8964 15379 8998 15413
rect 8964 15311 8998 15345
rect 8964 15243 8998 15277
rect 8964 15175 8998 15209
rect 8964 15107 8998 15141
rect 8964 15039 8998 15073
rect 8964 14971 8998 15005
rect 8964 14903 8998 14937
rect 9904 16254 9938 16288
rect 9904 16186 9938 16220
rect 9904 16118 9938 16152
rect 9904 16050 9938 16084
rect 11457 16310 11491 16344
rect 11457 16242 11491 16276
rect 11457 16174 11491 16208
rect 11457 16106 11491 16140
rect 17181 17604 17215 17638
rect 17181 17536 17215 17570
rect 17181 17468 17215 17502
rect 17181 17400 17215 17434
rect 17181 17332 17215 17366
rect 17181 17264 17215 17298
rect 17181 17196 17215 17230
rect 17181 17128 17215 17162
rect 17181 17060 17215 17094
rect 17181 16992 17215 17026
rect 17181 16924 17215 16958
rect 17181 16856 17215 16890
rect 17181 16788 17215 16822
rect 17181 16720 17215 16754
rect 17181 16652 17215 16686
rect 17181 16584 17215 16618
rect 17181 16516 17215 16550
rect 17181 16448 17215 16482
rect 17181 16380 17215 16414
rect 17181 16312 17215 16346
rect 17181 16244 17215 16278
rect 17181 16176 17215 16210
rect 17181 16082 17215 16142
rect 11491 16072 11581 16082
rect 11457 16048 11581 16072
rect 11615 16048 11649 16082
rect 11683 16048 11717 16082
rect 11751 16048 11785 16082
rect 11819 16048 11853 16082
rect 11887 16048 11921 16082
rect 11955 16048 11989 16082
rect 12023 16048 12057 16082
rect 12091 16048 12125 16082
rect 12159 16048 12193 16082
rect 12227 16048 12261 16082
rect 12295 16048 12329 16082
rect 12363 16048 12397 16082
rect 12431 16048 12465 16082
rect 12499 16048 12533 16082
rect 12567 16048 12601 16082
rect 12635 16048 12669 16082
rect 12703 16048 12737 16082
rect 12771 16048 12805 16082
rect 12839 16048 12873 16082
rect 12907 16048 12941 16082
rect 12975 16048 13009 16082
rect 13043 16048 13077 16082
rect 13111 16048 13145 16082
rect 13179 16048 13213 16082
rect 13247 16048 13281 16082
rect 13315 16048 13349 16082
rect 13383 16048 13417 16082
rect 13451 16048 13485 16082
rect 13519 16048 13553 16082
rect 13587 16048 13621 16082
rect 13655 16048 13689 16082
rect 13723 16048 13757 16082
rect 13791 16048 13825 16082
rect 13859 16048 13893 16082
rect 13927 16048 13961 16082
rect 13995 16048 14029 16082
rect 14063 16048 14097 16082
rect 14131 16048 14165 16082
rect 14199 16048 14233 16082
rect 14267 16048 14301 16082
rect 14335 16048 14369 16082
rect 14403 16048 14437 16082
rect 14471 16048 14505 16082
rect 14539 16048 14573 16082
rect 14607 16048 14641 16082
rect 14675 16048 14709 16082
rect 14743 16048 14777 16082
rect 14811 16048 14845 16082
rect 14879 16048 14913 16082
rect 14947 16048 14981 16082
rect 15015 16048 15049 16082
rect 15083 16048 15117 16082
rect 15151 16048 15185 16082
rect 15219 16048 15253 16082
rect 15287 16048 15321 16082
rect 15355 16048 15389 16082
rect 15423 16048 15457 16082
rect 15491 16048 15525 16082
rect 15559 16048 15593 16082
rect 15627 16048 15661 16082
rect 15695 16048 15729 16082
rect 15763 16048 15797 16082
rect 15831 16048 15865 16082
rect 15899 16048 15933 16082
rect 15967 16048 16001 16082
rect 16035 16048 16069 16082
rect 16103 16048 16137 16082
rect 16171 16048 16205 16082
rect 16239 16048 16273 16082
rect 16307 16048 16341 16082
rect 16375 16048 16409 16082
rect 16443 16048 16477 16082
rect 16511 16048 16545 16082
rect 16579 16048 16613 16082
rect 16647 16048 16681 16082
rect 16715 16048 16749 16082
rect 16783 16048 16817 16082
rect 16851 16048 16885 16082
rect 16919 16048 16953 16082
rect 16987 16048 17021 16082
rect 17055 16048 17089 16082
rect 17123 16048 17157 16082
rect 17191 16048 17215 16082
rect 17287 19236 17383 19260
rect 17321 19226 17383 19236
rect 17417 19226 17451 19260
rect 17485 19226 17519 19260
rect 17553 19226 17587 19260
rect 17621 19226 17655 19260
rect 17689 19226 17723 19260
rect 17757 19226 17791 19260
rect 17825 19226 17859 19260
rect 17893 19226 17927 19260
rect 17961 19226 17995 19260
rect 18029 19226 18063 19260
rect 18097 19226 18131 19260
rect 18165 19226 18199 19260
rect 18233 19226 18267 19260
rect 18301 19226 18335 19260
rect 18369 19226 18403 19260
rect 18437 19226 18471 19260
rect 18505 19226 18539 19260
rect 18573 19226 18607 19260
rect 18641 19226 18675 19260
rect 18709 19226 18743 19260
rect 18777 19226 18811 19260
rect 18845 19226 18879 19260
rect 18913 19226 18947 19260
rect 18981 19226 19015 19260
rect 19049 19226 19083 19260
rect 19117 19226 19151 19260
rect 19185 19226 19219 19260
rect 19253 19226 19287 19260
rect 19321 19226 19355 19260
rect 19389 19226 19423 19260
rect 19457 19226 19491 19260
rect 19525 19226 19559 19260
rect 19593 19226 19627 19260
rect 19661 19226 19695 19260
rect 19729 19226 19763 19260
rect 19797 19226 19831 19260
rect 19865 19226 19899 19260
rect 19933 19226 19967 19260
rect 20001 19226 20035 19260
rect 20069 19226 20103 19260
rect 20137 19226 20171 19260
rect 20205 19226 20229 19260
rect 17287 19168 17321 19202
rect 17287 19100 17321 19134
rect 17287 19032 17321 19066
rect 17287 18964 17321 18998
rect 17287 18896 17321 18930
rect 17287 18828 17321 18862
rect 17287 18760 17321 18794
rect 17287 18692 17321 18726
rect 17287 18624 17321 18658
rect 17287 18556 17321 18590
rect 17287 18488 17321 18522
rect 17287 18420 17321 18454
rect 17287 18352 17321 18386
rect 17287 18284 17321 18318
rect 17287 18216 17321 18250
rect 17287 18148 17321 18182
rect 17287 18080 17321 18114
rect 17287 18012 17321 18046
rect 17287 17944 17321 17978
rect 17287 17876 17321 17910
rect 17287 17808 17321 17842
rect 17287 17740 17321 17774
rect 17287 17672 17321 17706
rect 17287 17604 17321 17638
rect 17287 17536 17321 17570
rect 17287 17468 17321 17502
rect 17287 17400 17321 17434
rect 17287 17332 17321 17366
rect 17287 17264 17321 17298
rect 17287 17196 17321 17230
rect 17287 17128 17321 17162
rect 17287 17060 17321 17094
rect 17287 16992 17321 17026
rect 17287 16924 17321 16958
rect 17287 16856 17321 16890
rect 17287 16788 17321 16822
rect 17287 16720 17321 16754
rect 17287 16652 17321 16686
rect 17287 16584 17321 16618
rect 17287 16516 17321 16550
rect 17287 16448 17321 16482
rect 17287 16380 17321 16414
rect 17287 16312 17321 16346
rect 17287 16244 17321 16278
rect 17287 16176 17321 16210
rect 17287 16082 17321 16142
rect 20195 19140 20229 19226
rect 20195 19072 20229 19106
rect 20195 19004 20229 19038
rect 20195 18936 20229 18970
rect 20195 18868 20229 18902
rect 20195 18800 20229 18834
rect 20195 18732 20229 18766
rect 20195 18664 20229 18698
rect 20195 18596 20229 18630
rect 20195 18528 20229 18562
rect 20195 18460 20229 18494
rect 20195 18392 20229 18426
rect 20195 18324 20229 18358
rect 20195 18256 20229 18290
rect 20195 18188 20229 18222
rect 20195 18120 20229 18154
rect 20195 18052 20229 18086
rect 20195 17984 20229 18018
rect 20195 17916 20229 17950
rect 20195 17848 20229 17882
rect 20195 17780 20229 17814
rect 20195 17712 20229 17746
rect 20195 17602 20229 17678
rect 20195 17534 20229 17568
rect 20195 17466 20229 17500
rect 20195 17398 20229 17432
rect 20195 17330 20229 17364
rect 20195 17262 20229 17296
rect 20195 17194 20229 17228
rect 20195 17126 20229 17160
rect 20195 17058 20229 17092
rect 20195 16990 20229 17024
rect 20195 16922 20229 16956
rect 20195 16854 20229 16888
rect 20195 16786 20229 16820
rect 20195 16718 20229 16752
rect 20195 16650 20229 16684
rect 20195 16582 20229 16616
rect 20195 16514 20229 16548
rect 20195 16446 20229 16480
rect 20195 16378 20229 16412
rect 20195 16310 20229 16344
rect 20195 16242 20229 16276
rect 20195 16174 20229 16208
rect 20195 16106 20229 16140
rect 17287 16048 17311 16082
rect 17345 16048 17379 16082
rect 17413 16048 17447 16082
rect 17481 16048 17515 16082
rect 17549 16048 17583 16082
rect 17617 16048 17651 16082
rect 17685 16048 17719 16082
rect 17753 16048 17787 16082
rect 17821 16048 17855 16082
rect 17889 16048 17923 16082
rect 17957 16048 17991 16082
rect 18025 16048 18059 16082
rect 18093 16048 18127 16082
rect 18161 16048 18195 16082
rect 18229 16048 18263 16082
rect 18297 16048 18331 16082
rect 18365 16048 18399 16082
rect 18433 16048 18467 16082
rect 18501 16048 18535 16082
rect 18569 16048 18603 16082
rect 18637 16048 18671 16082
rect 18705 16048 18739 16082
rect 18773 16048 18807 16082
rect 18841 16048 18875 16082
rect 18909 16048 18943 16082
rect 18977 16048 19011 16082
rect 19045 16048 19079 16082
rect 19113 16048 19147 16082
rect 19181 16048 19215 16082
rect 19249 16048 19283 16082
rect 19317 16048 19351 16082
rect 19385 16048 19419 16082
rect 19453 16048 19487 16082
rect 19521 16048 19555 16082
rect 19589 16048 19623 16082
rect 19657 16048 19691 16082
rect 19725 16048 19759 16082
rect 19793 16048 19827 16082
rect 19861 16048 19895 16082
rect 19929 16048 19963 16082
rect 19997 16048 20031 16082
rect 20065 16048 20099 16082
rect 20133 16072 20195 16082
rect 20133 16048 20229 16072
rect 20301 19236 20374 19260
rect 20335 19226 20374 19236
rect 20408 19226 20442 19260
rect 20476 19226 20510 19260
rect 20544 19226 20578 19260
rect 20612 19226 20646 19260
rect 20680 19226 20714 19260
rect 20748 19226 20782 19260
rect 20816 19226 20850 19260
rect 20884 19226 20918 19260
rect 20952 19226 20986 19260
rect 21020 19226 21054 19260
rect 21088 19226 21122 19260
rect 21156 19226 21190 19260
rect 21224 19226 21258 19260
rect 21292 19226 21326 19260
rect 21360 19226 21394 19260
rect 21428 19226 21462 19260
rect 21496 19226 21530 19260
rect 21564 19226 21598 19260
rect 21632 19226 21666 19260
rect 21700 19226 21734 19260
rect 21768 19226 21802 19260
rect 21836 19226 21870 19260
rect 21904 19226 21938 19260
rect 21972 19226 22006 19260
rect 22040 19226 22074 19260
rect 22108 19226 22142 19260
rect 22176 19226 22210 19260
rect 22244 19226 22278 19260
rect 22312 19226 22346 19260
rect 22380 19226 22414 19260
rect 22448 19226 22482 19260
rect 22516 19226 22550 19260
rect 22584 19226 22618 19260
rect 22652 19226 22686 19260
rect 22720 19226 22754 19260
rect 22788 19226 22822 19260
rect 22856 19226 22890 19260
rect 22924 19226 22958 19260
rect 22992 19226 23026 19260
rect 23060 19226 23157 19260
rect 23191 19226 23225 19260
rect 23259 19226 23293 19260
rect 23327 19226 23361 19260
rect 23395 19226 23429 19260
rect 23463 19226 23497 19260
rect 23531 19226 23565 19260
rect 23599 19226 23633 19260
rect 23667 19226 23701 19260
rect 23735 19226 23769 19260
rect 23803 19226 23837 19260
rect 23871 19226 23905 19260
rect 23939 19226 23973 19260
rect 24007 19226 24041 19260
rect 24075 19226 24109 19260
rect 24143 19226 24177 19260
rect 24211 19226 24245 19260
rect 24279 19226 24313 19260
rect 24347 19226 24381 19260
rect 24415 19226 24449 19260
rect 24483 19226 24517 19260
rect 24551 19226 24585 19260
rect 24619 19226 24653 19260
rect 24687 19226 24721 19260
rect 24755 19226 24789 19260
rect 24823 19226 24857 19260
rect 24891 19226 24925 19260
rect 24959 19226 24993 19260
rect 25027 19226 25061 19260
rect 25095 19226 25129 19260
rect 25163 19226 25197 19260
rect 25231 19226 25265 19260
rect 25299 19226 25333 19260
rect 25367 19226 25401 19260
rect 25435 19226 25469 19260
rect 25503 19226 25537 19260
rect 25571 19226 25605 19260
rect 25639 19226 25673 19260
rect 25707 19226 25741 19260
rect 25775 19226 25809 19260
rect 25843 19226 25867 19260
rect 20301 19168 20335 19202
rect 20301 19100 20335 19134
rect 20301 19032 20335 19066
rect 20301 18964 20335 18998
rect 20301 18896 20335 18930
rect 20301 18828 20335 18862
rect 20301 18760 20335 18794
rect 20301 18692 20335 18726
rect 20301 18624 20335 18658
rect 20301 18556 20335 18590
rect 20301 18488 20335 18522
rect 20301 18420 20335 18454
rect 20301 18352 20335 18386
rect 20301 18284 20335 18318
rect 20301 18216 20335 18250
rect 20301 18148 20335 18182
rect 20301 18080 20335 18114
rect 20301 18012 20335 18046
rect 20301 17944 20335 17978
rect 20301 17876 20335 17910
rect 20301 17808 20335 17842
rect 20301 17740 20335 17774
rect 20301 17672 20335 17706
rect 20301 17604 20335 17638
rect 20301 17536 20335 17570
rect 20301 17468 20335 17502
rect 20301 17400 20335 17434
rect 20301 17332 20335 17366
rect 20301 17264 20335 17298
rect 20301 17196 20335 17230
rect 20301 17128 20335 17162
rect 20301 17060 20335 17094
rect 20301 16992 20335 17026
rect 20301 16924 20335 16958
rect 20301 16856 20335 16890
rect 20301 16788 20335 16822
rect 20301 16720 20335 16754
rect 20301 16652 20335 16686
rect 20301 16584 20335 16618
rect 20301 16516 20335 16550
rect 20301 16448 20335 16482
rect 20301 16380 20335 16414
rect 20301 16312 20335 16346
rect 20301 16244 20335 16278
rect 20301 16176 20335 16210
rect 20301 16082 20335 16142
rect 25833 19166 25867 19226
rect 25833 19098 25867 19132
rect 25833 19030 25867 19064
rect 25833 18962 25867 18996
rect 25833 18894 25867 18928
rect 25833 18826 25867 18860
rect 25833 18758 25867 18792
rect 25833 18690 25867 18724
rect 25833 18622 25867 18656
rect 25833 18554 25867 18588
rect 25833 18486 25867 18520
rect 25833 18418 25867 18452
rect 25833 18350 25867 18384
rect 25833 18282 25867 18316
rect 25833 18214 25867 18248
rect 25833 18146 25867 18180
rect 25833 18078 25867 18112
rect 25833 18010 25867 18044
rect 25833 17942 25867 17976
rect 25833 17874 25867 17908
rect 25833 17806 25867 17840
rect 25833 17738 25867 17772
rect 25833 17670 25867 17704
rect 25833 17602 25867 17636
rect 25833 17534 25867 17568
rect 25833 17466 25867 17500
rect 25833 17398 25867 17432
rect 25833 17330 25867 17364
rect 25833 17262 25867 17296
rect 25833 17194 25867 17228
rect 25833 17126 25867 17160
rect 25833 17058 25867 17092
rect 25833 16990 25867 17024
rect 25833 16922 25867 16956
rect 25833 16854 25867 16888
rect 25833 16786 25867 16820
rect 25833 16718 25867 16752
rect 25833 16650 25867 16684
rect 25833 16582 25867 16616
rect 25833 16514 25867 16548
rect 25833 16446 25867 16480
rect 25833 16378 25867 16412
rect 25833 16310 25867 16344
rect 25833 16242 25867 16276
rect 25833 16174 25867 16208
rect 25833 16106 25867 16140
rect 20301 16048 20325 16082
rect 20359 16048 20393 16082
rect 20427 16048 20461 16082
rect 20495 16048 20529 16082
rect 20563 16048 20597 16082
rect 20631 16048 20665 16082
rect 20699 16048 20733 16082
rect 20767 16048 20801 16082
rect 20835 16048 20869 16082
rect 20903 16048 20937 16082
rect 20971 16048 21005 16082
rect 21039 16048 21073 16082
rect 21107 16048 21141 16082
rect 21175 16048 21209 16082
rect 21243 16048 21277 16082
rect 21311 16048 21345 16082
rect 21379 16048 21413 16082
rect 21447 16048 21481 16082
rect 21515 16048 21549 16082
rect 21583 16048 21617 16082
rect 21651 16048 21685 16082
rect 21719 16048 21753 16082
rect 21787 16048 21821 16082
rect 21855 16048 21889 16082
rect 21923 16048 21957 16082
rect 21991 16048 22025 16082
rect 22059 16048 22093 16082
rect 22127 16048 22161 16082
rect 22195 16048 22229 16082
rect 22263 16048 22297 16082
rect 22331 16048 22365 16082
rect 22399 16048 22433 16082
rect 22467 16048 22501 16082
rect 22535 16048 22569 16082
rect 22603 16048 22637 16082
rect 22671 16048 22705 16082
rect 22739 16048 22773 16082
rect 22807 16048 22841 16082
rect 22875 16048 22909 16082
rect 22943 16048 22977 16082
rect 23011 16048 23045 16082
rect 23079 16048 23113 16082
rect 23147 16048 23181 16082
rect 23215 16048 23249 16082
rect 23283 16048 23317 16082
rect 23351 16048 23385 16082
rect 23419 16048 23453 16082
rect 23487 16048 23521 16082
rect 23555 16048 23589 16082
rect 23623 16048 23657 16082
rect 23691 16048 23725 16082
rect 23759 16048 23793 16082
rect 23827 16048 23861 16082
rect 23895 16048 23929 16082
rect 23963 16048 23997 16082
rect 24031 16048 24065 16082
rect 24099 16048 24133 16082
rect 24167 16048 24201 16082
rect 24235 16048 24269 16082
rect 24303 16048 24337 16082
rect 24371 16048 24405 16082
rect 24439 16048 24473 16082
rect 24507 16048 24541 16082
rect 24575 16048 24609 16082
rect 24643 16048 24677 16082
rect 24711 16048 24745 16082
rect 24779 16048 24813 16082
rect 24847 16048 24881 16082
rect 24915 16048 24949 16082
rect 24983 16048 25017 16082
rect 25051 16048 25085 16082
rect 25119 16048 25153 16082
rect 25187 16048 25221 16082
rect 25255 16048 25289 16082
rect 25323 16048 25357 16082
rect 25391 16048 25425 16082
rect 25459 16048 25493 16082
rect 25527 16048 25561 16082
rect 25595 16048 25629 16082
rect 25663 16048 25697 16082
rect 25731 16048 25765 16082
rect 25799 16072 25833 16082
rect 25799 16048 25867 16072
rect 9904 15982 9938 16016
rect 9904 15914 9938 15948
rect 9904 15846 9938 15880
rect 9904 15778 9938 15812
rect 9904 15710 9938 15744
rect 9904 15642 9938 15676
rect 9904 15574 9938 15608
rect 9904 15506 9938 15540
rect 9904 15438 9938 15472
rect 9904 15370 9938 15404
rect 9904 15302 9938 15336
rect 11457 15942 11481 15976
rect 11515 15942 11549 15976
rect 11583 15942 11617 15976
rect 11651 15942 11685 15976
rect 11719 15942 11753 15976
rect 11787 15942 11821 15976
rect 11855 15942 11889 15976
rect 11923 15942 11957 15976
rect 11991 15942 12025 15976
rect 12059 15942 12093 15976
rect 12127 15942 12161 15976
rect 12195 15942 12229 15976
rect 12263 15942 12297 15976
rect 12331 15942 12365 15976
rect 12399 15942 12433 15976
rect 12467 15942 12501 15976
rect 12535 15942 12649 15976
rect 12683 15942 12717 15976
rect 12751 15942 12785 15976
rect 12819 15942 12853 15976
rect 12887 15942 12921 15976
rect 12955 15942 12989 15976
rect 13023 15942 13057 15976
rect 13091 15942 13125 15976
rect 13159 15942 13193 15976
rect 13227 15942 13261 15976
rect 13295 15942 13329 15976
rect 13363 15942 13397 15976
rect 13431 15942 13465 15976
rect 13499 15942 13533 15976
rect 13567 15942 13601 15976
rect 13635 15942 13669 15976
rect 13703 15952 13793 15976
rect 17215 15975 17239 15976
rect 13703 15942 13759 15952
rect 11457 15902 11491 15942
rect 11457 15834 11491 15868
rect 11457 15766 11491 15800
rect 11457 15698 11491 15732
rect 11457 15630 11491 15664
rect 11457 15562 11491 15596
rect 11457 15494 11491 15528
rect 11457 15426 11491 15460
rect 11457 15358 11491 15392
rect 11457 15290 11491 15324
rect 9904 15234 9938 15268
rect 11457 15222 11491 15256
rect 9904 15166 9938 15200
rect 9904 15098 9938 15132
rect 11457 15154 11491 15188
rect 11457 15086 11491 15120
rect 9904 15030 9938 15064
rect 9904 14962 9938 14996
rect 9904 14879 9938 14928
rect 8998 14869 9064 14879
rect 8964 14845 9064 14869
rect 9098 14845 9132 14879
rect 9166 14845 9200 14879
rect 9234 14845 9268 14879
rect 9302 14845 9336 14879
rect 9370 14845 9404 14879
rect 9438 14845 9472 14879
rect 9506 14845 9540 14879
rect 9574 14845 9608 14879
rect 9642 14845 9676 14879
rect 9710 14845 9744 14879
rect 9778 14845 9812 14879
rect 9846 14845 9880 14879
rect 9914 14845 9938 14879
rect 11457 15018 11491 15052
rect 11457 14950 11491 14984
rect 11457 14882 11491 14916
rect 13759 15884 13793 15918
rect 13759 15816 13793 15850
rect 13759 15748 13793 15782
rect 13759 15680 13793 15714
rect 13759 15612 13793 15646
rect 13759 15544 13793 15578
rect 13759 15476 13793 15510
rect 13759 15408 13793 15442
rect 13759 15340 13793 15374
rect 13759 15272 13793 15306
rect 13759 15204 13793 15238
rect 13759 15136 13793 15170
rect 13759 15068 13793 15102
rect 13759 15000 13793 15034
rect 13759 14932 13793 14966
rect 13759 14858 13793 14898
rect 11491 14848 11559 14858
rect 11457 14824 11559 14848
rect 11593 14824 11627 14858
rect 11661 14824 11695 14858
rect 11729 14824 11763 14858
rect 11797 14824 11831 14858
rect 11865 14824 11899 14858
rect 11933 14824 11967 14858
rect 12001 14824 12035 14858
rect 12069 14824 12103 14858
rect 12137 14824 12171 14858
rect 12205 14824 12239 14858
rect 12273 14824 12307 14858
rect 12341 14824 12375 14858
rect 12409 14824 12443 14858
rect 12477 14824 12511 14858
rect 12545 14824 12579 14858
rect 12613 14824 12647 14858
rect 12681 14824 12715 14858
rect 12749 14824 12783 14858
rect 12817 14824 12851 14858
rect 12885 14824 12919 14858
rect 12953 14824 12987 14858
rect 13021 14824 13055 14858
rect 13089 14824 13123 14858
rect 13157 14824 13191 14858
rect 13225 14824 13259 14858
rect 13293 14824 13327 14858
rect 13361 14824 13395 14858
rect 13429 14824 13463 14858
rect 13497 14824 13531 14858
rect 13565 14824 13599 14858
rect 13633 14824 13667 14858
rect 13701 14824 13735 14858
rect 13769 14824 13793 14858
rect 13865 15940 13889 15974
rect 13923 15940 13957 15974
rect 13991 15940 14025 15974
rect 14059 15940 14093 15974
rect 14127 15940 14161 15974
rect 14195 15940 14229 15974
rect 14263 15940 14297 15974
rect 14331 15940 14365 15974
rect 14399 15940 14433 15974
rect 14467 15940 14501 15974
rect 14535 15940 14569 15974
rect 14603 15940 14637 15974
rect 14671 15940 14705 15974
rect 14739 15940 14773 15974
rect 14807 15950 14931 15974
rect 14807 15940 14897 15950
rect 13865 15865 13899 15940
rect 13865 15797 13899 15831
rect 13865 15729 13899 15763
rect 13865 15661 13899 15695
rect 13865 15593 13899 15627
rect 13865 15525 13899 15559
rect 13865 15457 13899 15491
rect 13865 15358 13899 15423
rect 13865 15290 13899 15324
rect 13865 15222 13899 15256
rect 13865 15154 13899 15188
rect 13865 15086 13899 15120
rect 13865 15018 13899 15052
rect 13865 14950 13899 14984
rect 13865 14882 13899 14916
rect 14897 15882 14931 15916
rect 14897 15814 14931 15848
rect 14897 15746 14931 15780
rect 14897 15678 14931 15712
rect 14897 15610 14931 15644
rect 14897 15542 14931 15576
rect 14897 15474 14931 15508
rect 14897 15406 14931 15440
rect 14897 15338 14931 15372
rect 14897 15270 14931 15304
rect 14897 15202 14931 15236
rect 14897 15134 14931 15168
rect 14897 15066 14931 15100
rect 14897 14998 14931 15032
rect 14897 14930 14931 14964
rect 14897 14858 14931 14896
rect 13899 14848 13989 14858
rect 13865 14824 13989 14848
rect 14023 14824 14057 14858
rect 14091 14824 14125 14858
rect 14159 14824 14193 14858
rect 14227 14824 14261 14858
rect 14295 14824 14329 14858
rect 14363 14824 14397 14858
rect 14431 14824 14465 14858
rect 14499 14824 14533 14858
rect 14567 14824 14601 14858
rect 14635 14824 14669 14858
rect 14703 14824 14737 14858
rect 14771 14824 14805 14858
rect 14839 14824 14873 14858
rect 14907 14824 14931 14858
rect 15003 15941 15027 15975
rect 15061 15941 15095 15975
rect 15129 15941 15163 15975
rect 15197 15941 15231 15975
rect 15265 15941 15299 15975
rect 15333 15941 15367 15975
rect 15401 15941 15435 15975
rect 15469 15941 15503 15975
rect 15537 15941 15571 15975
rect 15605 15941 15639 15975
rect 15673 15941 15707 15975
rect 15741 15941 15775 15975
rect 15809 15941 15843 15975
rect 15877 15941 15911 15975
rect 15945 15941 15979 15975
rect 16013 15941 16047 15975
rect 16081 15941 16115 15975
rect 16149 15941 16183 15975
rect 16217 15941 16251 15975
rect 16285 15941 16319 15975
rect 16353 15941 16387 15975
rect 16421 15941 16455 15975
rect 16489 15941 16523 15975
rect 16557 15941 16591 15975
rect 16625 15941 16659 15975
rect 16693 15941 16727 15975
rect 16761 15941 16795 15975
rect 16829 15941 16863 15975
rect 16897 15941 16931 15975
rect 16965 15941 16999 15975
rect 17033 15941 17067 15975
rect 17101 15941 17135 15975
rect 17169 15942 17239 15975
rect 17273 15942 17307 15976
rect 17341 15942 17375 15976
rect 17409 15942 17443 15976
rect 17477 15942 17511 15976
rect 17545 15942 17579 15976
rect 17613 15942 17647 15976
rect 17681 15942 17715 15976
rect 17749 15942 17783 15976
rect 17817 15942 17851 15976
rect 17885 15942 17919 15976
rect 17953 15942 17987 15976
rect 18021 15942 18055 15976
rect 18089 15952 18205 15976
rect 18089 15942 18171 15952
rect 17169 15941 17249 15942
rect 15003 15902 15037 15941
rect 15003 15834 15037 15868
rect 15003 15766 15037 15800
rect 15003 15698 15037 15732
rect 15003 15630 15037 15664
rect 15003 15562 15037 15596
rect 15003 15494 15037 15528
rect 15003 15426 15037 15460
rect 15003 15358 15037 15392
rect 15003 15290 15037 15324
rect 15003 15222 15037 15256
rect 15003 15154 15037 15188
rect 15003 15086 15037 15120
rect 15003 15018 15037 15052
rect 15003 14950 15037 14984
rect 15003 14882 15037 14916
rect 18171 15884 18205 15918
rect 18171 15816 18205 15850
rect 18171 15748 18205 15782
rect 18171 15680 18205 15714
rect 18171 15612 18205 15646
rect 18171 15544 18205 15578
rect 18171 15476 18205 15510
rect 18171 15408 18205 15442
rect 18171 15340 18205 15374
rect 18171 15272 18205 15306
rect 18171 15204 18205 15238
rect 18171 15136 18205 15170
rect 18171 15068 18205 15102
rect 18171 15000 18205 15034
rect 18171 14932 18205 14966
rect 18171 14858 18205 14898
rect 15037 14848 15118 14858
rect 15003 14824 15118 14848
rect 15152 14824 15186 14858
rect 15220 14824 15254 14858
rect 15288 14824 15322 14858
rect 15356 14824 15390 14858
rect 15424 14824 15458 14858
rect 15492 14824 15526 14858
rect 15560 14824 15594 14858
rect 15628 14824 15662 14858
rect 15696 14824 15730 14858
rect 15764 14824 15798 14858
rect 15832 14824 15866 14858
rect 15900 14824 15934 14858
rect 15968 14824 16002 14858
rect 16036 14824 16070 14858
rect 16104 14824 16138 14858
rect 16172 14824 16206 14858
rect 16240 14824 16274 14858
rect 16308 14824 16342 14858
rect 16376 14824 16410 14858
rect 16444 14824 16478 14858
rect 16512 14824 16546 14858
rect 16580 14824 16651 14858
rect 16685 14824 16719 14858
rect 16753 14824 16787 14858
rect 16821 14824 16855 14858
rect 16889 14824 16923 14858
rect 16957 14824 16991 14858
rect 17025 14824 17059 14858
rect 17093 14824 17127 14858
rect 17161 14824 17195 14858
rect 17229 14824 17263 14858
rect 17297 14824 17331 14858
rect 17365 14824 17399 14858
rect 17433 14824 17467 14858
rect 17501 14824 17535 14858
rect 17569 14824 17603 14858
rect 17637 14824 17671 14858
rect 17705 14824 17739 14858
rect 17773 14824 17807 14858
rect 17841 14824 17875 14858
rect 17909 14824 17943 14858
rect 17977 14824 18011 14858
rect 18045 14824 18079 14858
rect 18113 14824 18147 14858
rect 18181 14824 18205 14858
<< psubdiffcont >>
rect 6976 33058 7010 33092
rect 7044 33058 7078 33092
rect 7112 33058 7146 33092
rect 7180 33058 7214 33092
rect 7248 33058 7282 33092
rect 7316 33058 7350 33092
rect 7384 33058 7418 33092
rect 7452 33058 7486 33092
rect 7520 33058 7554 33092
rect 7662 33064 7696 33098
rect 7730 33064 7764 33098
rect 7798 33064 7832 33098
rect 7914 33058 7948 33092
rect 6952 32942 6986 32976
rect 8038 32982 8072 33016
rect 6952 32874 6986 32908
rect 6952 32806 6986 32840
rect 6952 32738 6986 32772
rect 6952 32670 6986 32704
rect 6952 32602 6986 32636
rect 6952 32534 6986 32568
rect 6952 32466 6986 32500
rect 6952 32398 6986 32432
rect 6952 32330 6986 32364
rect 6952 32262 6986 32296
rect 6952 32194 6986 32228
rect 6952 32126 6986 32160
rect 6952 32058 6986 32092
rect 6952 31990 6986 32024
rect 6878 31898 6912 31932
rect 6952 31922 6986 31956
rect 8038 32914 8072 32948
rect 8038 32846 8072 32880
rect 9458 33004 9492 33038
rect 9526 33004 9560 33038
rect 9594 33004 9628 33038
rect 9662 33004 9696 33038
rect 9730 33004 9764 33038
rect 9798 33004 9832 33038
rect 9866 33004 9900 33038
rect 9934 33004 9968 33038
rect 10002 33004 10036 33038
rect 10070 33004 10104 33038
rect 10138 33004 10172 33038
rect 10206 33004 10240 33038
rect 10274 33004 10308 33038
rect 10342 33004 10376 33038
rect 10410 33004 10444 33038
rect 10478 33004 10512 33038
rect 10546 33004 10580 33038
rect 10614 33004 10648 33038
rect 10682 33004 10716 33038
rect 10750 33004 10784 33038
rect 10818 33004 10852 33038
rect 10886 33004 10920 33038
rect 10954 33004 10988 33038
rect 11022 33004 11056 33038
rect 11090 33004 11124 33038
rect 11158 33004 11192 33038
rect 9434 32893 9468 32927
rect 11242 32980 11276 33014
rect 8038 32778 8072 32812
rect 8038 32710 8072 32744
rect 9650 32876 9684 32910
rect 9718 32876 9752 32910
rect 9786 32876 9820 32910
rect 9854 32876 9888 32910
rect 9922 32876 9956 32910
rect 10044 32876 10078 32910
rect 10112 32876 10146 32910
rect 10180 32876 10214 32910
rect 10248 32876 10282 32910
rect 10400 32876 10434 32910
rect 10468 32876 10502 32910
rect 10536 32876 10570 32910
rect 10604 32876 10638 32910
rect 10743 32876 10777 32910
rect 10811 32876 10845 32910
rect 10879 32876 10913 32910
rect 10947 32876 10981 32910
rect 11015 32876 11049 32910
rect 11242 32912 11276 32946
rect 9434 32825 9468 32859
rect 11242 32844 11276 32878
rect 9434 32757 9468 32791
rect 8038 32642 8072 32676
rect 9434 32689 9468 32723
rect 8038 32574 8072 32608
rect 8038 32506 8072 32540
rect 8038 32438 8072 32472
rect 8038 32370 8072 32404
rect 8038 32302 8072 32336
rect 8038 32234 8072 32268
rect 8038 32166 8072 32200
rect 8038 32098 8072 32132
rect 8038 32030 8072 32064
rect 8038 31929 8072 31963
rect 6854 31793 6888 31827
rect 6854 31725 6888 31759
rect 6854 31657 6888 31691
rect 6854 31589 6888 31623
rect 8038 31861 8072 31895
rect 8038 31793 8072 31827
rect 8038 31725 8072 31759
rect 8038 31657 8072 31691
rect 6928 31565 6962 31599
rect 6996 31565 7030 31599
rect 7064 31565 7098 31599
rect 7132 31565 7166 31599
rect 7200 31565 7234 31599
rect 7268 31565 7302 31599
rect 7336 31565 7370 31599
rect 7360 31434 7394 31468
rect 7360 31366 7394 31400
rect 7360 31298 7394 31332
rect 7360 31230 7394 31264
rect 7360 31162 7394 31196
rect 7360 31094 7394 31128
rect 7360 31026 7394 31060
rect 7360 30958 7394 30992
rect 8038 31589 8072 31623
rect 8038 31521 8072 31555
rect 8038 31453 8072 31487
rect 8038 31385 8072 31419
rect 8038 31317 8072 31351
rect 8038 31249 8072 31283
rect 8038 31181 8072 31215
rect 8038 31113 8072 31147
rect 8038 31045 8072 31079
rect 9434 32621 9468 32655
rect 9434 32553 9468 32587
rect 9434 32485 9468 32519
rect 9434 32417 9468 32451
rect 9434 32349 9468 32383
rect 9434 32281 9468 32315
rect 9434 32213 9468 32247
rect 9434 32145 9468 32179
rect 9434 32077 9468 32111
rect 9434 32009 9468 32043
rect 9434 31941 9468 31975
rect 9434 31873 9468 31907
rect 9434 31805 9468 31839
rect 9434 31737 9468 31771
rect 9434 31669 9468 31703
rect 9434 31601 9468 31635
rect 9434 31533 9468 31567
rect 9434 31465 9468 31499
rect 9434 31397 9468 31431
rect 11242 32776 11276 32810
rect 11242 32708 11276 32742
rect 11242 32640 11276 32674
rect 11242 32572 11276 32606
rect 11242 32504 11276 32538
rect 11242 32436 11276 32470
rect 11242 32368 11276 32402
rect 11242 32300 11276 32334
rect 11242 32232 11276 32266
rect 11242 32164 11276 32198
rect 11242 32096 11276 32130
rect 11242 32028 11276 32062
rect 11242 31960 11276 31994
rect 11242 31892 11276 31926
rect 11242 31824 11276 31858
rect 11242 31756 11276 31790
rect 11242 31688 11276 31722
rect 11242 31620 11276 31654
rect 11242 31552 11276 31586
rect 11330 32980 11364 33014
rect 11422 33004 11456 33038
rect 11490 33004 11524 33038
rect 11558 33004 11592 33038
rect 11626 33004 11660 33038
rect 11694 33004 11728 33038
rect 11762 33004 11796 33038
rect 11830 33004 11864 33038
rect 11898 33004 11932 33038
rect 11966 33004 12000 33038
rect 12034 33004 12068 33038
rect 12102 33004 12136 33038
rect 12170 33004 12204 33038
rect 12238 33004 12272 33038
rect 12306 33004 12340 33038
rect 12374 33004 12408 33038
rect 12442 33004 12476 33038
rect 12510 33004 12544 33038
rect 12578 33004 12612 33038
rect 12646 33004 12680 33038
rect 12714 33004 12748 33038
rect 12782 33004 12816 33038
rect 12850 33004 12884 33038
rect 12918 33004 12952 33038
rect 12986 33004 13020 33038
rect 13054 33004 13088 33038
rect 13122 33004 13156 33038
rect 13190 33004 13224 33038
rect 13258 33004 13292 33038
rect 13326 33004 13360 33038
rect 13394 33004 13428 33038
rect 13462 33004 13496 33038
rect 13530 33004 13564 33038
rect 13598 33004 13632 33038
rect 13666 33004 13700 33038
rect 13734 33004 13768 33038
rect 13802 33004 13836 33038
rect 13870 33004 13904 33038
rect 13938 33004 13972 33038
rect 14006 33004 14040 33038
rect 14074 33004 14108 33038
rect 14142 33004 14176 33038
rect 14210 33004 14244 33038
rect 14278 33004 14312 33038
rect 14346 33004 14380 33038
rect 14414 33004 14448 33038
rect 14482 33004 14516 33038
rect 14550 33004 14584 33038
rect 14618 33004 14652 33038
rect 14686 33004 14720 33038
rect 14754 33004 14788 33038
rect 14822 33004 14856 33038
rect 14890 33004 14924 33038
rect 14958 33004 14992 33038
rect 15026 33004 15060 33038
rect 15094 33004 15128 33038
rect 15162 33004 15196 33038
rect 15230 33004 15264 33038
rect 15298 33004 15332 33038
rect 15366 33004 15400 33038
rect 15434 33004 15468 33038
rect 15502 33004 15536 33038
rect 15570 33004 15604 33038
rect 15638 33004 15672 33038
rect 15706 33004 15740 33038
rect 15774 33004 15808 33038
rect 15842 33004 15876 33038
rect 15910 33004 15944 33038
rect 15978 33004 16012 33038
rect 16046 33004 16080 33038
rect 16114 33004 16148 33038
rect 16182 33004 16216 33038
rect 16250 33004 16284 33038
rect 16318 33004 16352 33038
rect 11330 32912 11364 32946
rect 11330 32844 11364 32878
rect 16342 32936 16376 32970
rect 16342 32868 16376 32902
rect 11330 32776 11364 32810
rect 11330 32708 11364 32742
rect 11330 32640 11364 32674
rect 11330 32572 11364 32606
rect 11330 32504 11364 32538
rect 11330 32436 11364 32470
rect 11330 32368 11364 32402
rect 16342 32800 16376 32834
rect 16342 32732 16376 32766
rect 16342 32664 16376 32698
rect 16342 32596 16376 32630
rect 16342 32528 16376 32562
rect 16342 32460 16376 32494
rect 16342 32392 16376 32426
rect 11330 32300 11364 32334
rect 16342 32324 16376 32358
rect 11330 32232 11364 32266
rect 11330 32164 11364 32198
rect 11330 32096 11364 32130
rect 11330 32028 11364 32062
rect 11330 31960 11364 31994
rect 11330 31892 11364 31926
rect 11330 31824 11364 31858
rect 16342 32256 16376 32290
rect 16342 32188 16376 32222
rect 16342 32120 16376 32154
rect 16342 32052 16376 32086
rect 16342 31984 16376 32018
rect 16342 31916 16376 31950
rect 16342 31848 16376 31882
rect 11330 31756 11364 31790
rect 16342 31780 16376 31814
rect 11330 31688 11364 31722
rect 11469 31678 11503 31712
rect 11537 31678 11571 31712
rect 11605 31678 11639 31712
rect 11673 31678 11707 31712
rect 11741 31678 11775 31712
rect 11809 31678 11843 31712
rect 11877 31678 11911 31712
rect 11945 31678 11979 31712
rect 12063 31678 12097 31712
rect 12131 31678 12165 31712
rect 12199 31678 12233 31712
rect 12267 31678 12301 31712
rect 12335 31678 12369 31712
rect 12403 31678 12437 31712
rect 12471 31678 12505 31712
rect 12606 31678 12640 31712
rect 12674 31678 12708 31712
rect 12742 31678 12776 31712
rect 12810 31678 12844 31712
rect 12878 31678 12912 31712
rect 12946 31678 12980 31712
rect 13014 31678 13048 31712
rect 13082 31678 13116 31712
rect 13260 31678 13294 31712
rect 13328 31678 13362 31712
rect 13396 31678 13430 31712
rect 13464 31678 13498 31712
rect 13532 31678 13566 31712
rect 13600 31678 13634 31712
rect 13668 31678 13702 31712
rect 13736 31678 13770 31712
rect 13841 31678 13875 31712
rect 13909 31678 13943 31712
rect 13977 31678 14011 31712
rect 14045 31678 14079 31712
rect 14113 31678 14147 31712
rect 14181 31678 14215 31712
rect 14249 31678 14283 31712
rect 14317 31678 14351 31712
rect 16342 31712 16376 31746
rect 11330 31620 11364 31654
rect 16342 31644 16376 31678
rect 11354 31552 11388 31586
rect 11422 31552 11456 31586
rect 11490 31552 11524 31586
rect 11558 31552 11592 31586
rect 11626 31552 11660 31586
rect 11694 31552 11728 31586
rect 11762 31552 11796 31586
rect 11830 31552 11864 31586
rect 11898 31552 11932 31586
rect 11966 31552 12000 31586
rect 12034 31552 12068 31586
rect 12102 31552 12136 31586
rect 12170 31552 12204 31586
rect 12238 31552 12272 31586
rect 12306 31552 12340 31586
rect 12374 31552 12408 31586
rect 12442 31552 12476 31586
rect 12510 31552 12544 31586
rect 12578 31552 12612 31586
rect 12646 31552 12680 31586
rect 12714 31552 12748 31586
rect 12782 31552 12816 31586
rect 12850 31552 12884 31586
rect 12918 31552 12952 31586
rect 12986 31552 13020 31586
rect 13054 31552 13088 31586
rect 13122 31552 13156 31586
rect 13190 31552 13224 31586
rect 13258 31552 13292 31586
rect 13326 31552 13360 31586
rect 13394 31552 13428 31586
rect 13462 31552 13496 31586
rect 13530 31552 13564 31586
rect 13598 31552 13632 31586
rect 13666 31552 13700 31586
rect 13734 31552 13768 31586
rect 13877 31552 13911 31586
rect 13945 31552 13979 31586
rect 14013 31552 14047 31586
rect 14081 31552 14115 31586
rect 14149 31552 14183 31586
rect 14217 31552 14251 31586
rect 14285 31552 14319 31586
rect 14353 31552 14387 31586
rect 14421 31552 14455 31586
rect 14489 31552 14523 31586
rect 14557 31552 14591 31586
rect 14625 31552 14659 31586
rect 14693 31552 14727 31586
rect 14761 31552 14795 31586
rect 14829 31552 14863 31586
rect 14897 31552 14931 31586
rect 14965 31552 14999 31586
rect 15033 31552 15067 31586
rect 15101 31552 15135 31586
rect 15169 31552 15203 31586
rect 15237 31552 15271 31586
rect 15305 31552 15339 31586
rect 15373 31552 15407 31586
rect 15441 31552 15475 31586
rect 15509 31552 15543 31586
rect 15577 31552 15611 31586
rect 15645 31552 15679 31586
rect 15713 31552 15747 31586
rect 15781 31552 15815 31586
rect 15849 31552 15883 31586
rect 15917 31552 15951 31586
rect 15985 31552 16019 31586
rect 16053 31552 16087 31586
rect 16121 31552 16155 31586
rect 16189 31552 16223 31586
rect 16257 31552 16291 31586
rect 16342 31576 16376 31610
rect 11242 31484 11276 31518
rect 11242 31416 11276 31450
rect 9434 31329 9468 31363
rect 11242 31348 11276 31382
rect 9434 31261 9468 31295
rect 9434 31160 9468 31194
rect 11242 31280 11276 31314
rect 11242 31212 11276 31246
rect 12777 31346 12811 31380
rect 12845 31346 12879 31380
rect 12913 31346 12947 31380
rect 12981 31346 13015 31380
rect 13049 31346 13083 31380
rect 13117 31346 13151 31380
rect 13185 31346 13219 31380
rect 13253 31346 13287 31380
rect 13321 31346 13355 31380
rect 13389 31346 13423 31380
rect 13457 31346 13491 31380
rect 13525 31346 13559 31380
rect 13593 31346 13627 31380
rect 13661 31346 13695 31380
rect 13729 31346 13763 31380
rect 13797 31346 13831 31380
rect 13865 31346 13899 31380
rect 13933 31346 13967 31380
rect 14001 31346 14035 31380
rect 14069 31346 14103 31380
rect 14137 31346 14171 31380
rect 14205 31346 14239 31380
rect 14273 31346 14307 31380
rect 14341 31346 14375 31380
rect 14409 31346 14443 31380
rect 14477 31346 14511 31380
rect 12668 31232 12702 31266
rect 9434 31092 9468 31126
rect 11242 31144 11276 31178
rect 12668 31164 12702 31198
rect 14586 31232 14620 31266
rect 9434 31024 9468 31058
rect 7331 30809 7365 30843
rect 7331 30741 7365 30775
rect 7331 30673 7365 30707
rect 8067 30910 8101 30944
rect 8067 30842 8101 30876
rect 8067 30774 8101 30808
rect 7431 30649 7465 30683
rect 7499 30649 7533 30683
rect 7567 30649 7601 30683
rect 7635 30649 7669 30683
rect 7703 30649 7737 30683
rect 7771 30649 7805 30683
rect 7839 30649 7873 30683
rect 7907 30649 7941 30683
rect 7975 30649 8009 30683
rect 8043 30649 8077 30683
rect 9434 30956 9468 30990
rect 9434 30888 9468 30922
rect 9434 30820 9468 30854
rect 9434 30752 9468 30786
rect 9434 30684 9468 30718
rect 9434 30616 9468 30650
rect 9434 30548 9468 30582
rect 9434 30480 9468 30514
rect 9434 30412 9468 30446
rect 9434 30344 9468 30378
rect 9434 30276 9468 30310
rect 9434 30208 9468 30242
rect 9434 30140 9468 30174
rect 9434 30072 9468 30106
rect 9434 30004 9468 30038
rect 9434 29936 9468 29970
rect 9434 29868 9468 29902
rect 9434 29800 9468 29834
rect 9434 29732 9468 29766
rect 9434 29664 9468 29698
rect 11242 31076 11276 31110
rect 14586 31164 14620 31198
rect 12777 31050 12811 31084
rect 12845 31050 12879 31084
rect 12913 31050 12947 31084
rect 12981 31050 13015 31084
rect 13049 31050 13083 31084
rect 13117 31050 13151 31084
rect 13185 31050 13219 31084
rect 13253 31050 13287 31084
rect 13321 31050 13355 31084
rect 13389 31050 13423 31084
rect 13457 31050 13491 31084
rect 13525 31050 13559 31084
rect 13593 31050 13627 31084
rect 13661 31050 13695 31084
rect 13729 31050 13763 31084
rect 13797 31050 13831 31084
rect 13865 31050 13899 31084
rect 13933 31050 13967 31084
rect 14001 31050 14035 31084
rect 14069 31050 14103 31084
rect 14137 31050 14171 31084
rect 14205 31050 14239 31084
rect 14273 31050 14307 31084
rect 14341 31050 14375 31084
rect 14409 31050 14443 31084
rect 14477 31050 14511 31084
rect 11242 31008 11276 31042
rect 11242 30940 11276 30974
rect 11242 30872 11276 30906
rect 11242 30804 11276 30838
rect 11242 30736 11276 30770
rect 11242 30668 11276 30702
rect 11242 30600 11276 30634
rect 11242 30532 11276 30566
rect 11242 30464 11276 30498
rect 11242 30396 11276 30430
rect 11242 30328 11276 30362
rect 11242 30260 11276 30294
rect 11242 30192 11276 30226
rect 11242 30124 11276 30158
rect 11242 30056 11276 30090
rect 11242 29988 11276 30022
rect 11242 29920 11276 29954
rect 11242 29852 11276 29886
rect 11242 29784 11276 29818
rect 11242 29716 11276 29750
rect 9434 29596 9468 29630
rect 11242 29648 11276 29682
rect 9434 29528 9468 29562
rect 9667 29564 9701 29598
rect 9735 29564 9769 29598
rect 9803 29564 9837 29598
rect 9871 29564 9905 29598
rect 9939 29564 9973 29598
rect 10078 29564 10112 29598
rect 10146 29564 10180 29598
rect 10214 29564 10248 29598
rect 10282 29564 10316 29598
rect 10417 29564 10451 29598
rect 10485 29564 10519 29598
rect 10553 29564 10587 29598
rect 10621 29564 10655 29598
rect 10743 29564 10777 29598
rect 10811 29564 10845 29598
rect 10879 29564 10913 29598
rect 10947 29564 10981 29598
rect 11015 29564 11049 29598
rect 11242 29580 11276 29614
rect 9434 29460 9468 29494
rect 11242 29512 11276 29546
rect 9518 29436 9552 29470
rect 9586 29436 9620 29470
rect 9654 29436 9688 29470
rect 9722 29436 9756 29470
rect 9790 29436 9824 29470
rect 9858 29436 9892 29470
rect 9926 29436 9960 29470
rect 9994 29436 10028 29470
rect 10062 29436 10096 29470
rect 10130 29436 10164 29470
rect 10198 29436 10232 29470
rect 10266 29436 10300 29470
rect 10334 29436 10368 29470
rect 10402 29436 10436 29470
rect 10470 29436 10504 29470
rect 10538 29436 10572 29470
rect 10606 29436 10640 29470
rect 10674 29436 10708 29470
rect 10742 29436 10776 29470
rect 10810 29436 10844 29470
rect 10878 29436 10912 29470
rect 10946 29436 10980 29470
rect 11014 29436 11048 29470
rect 11082 29436 11116 29470
rect 11150 29436 11184 29470
rect 11218 29436 11252 29470
rect 8988 14682 9022 14716
rect 9056 14682 9090 14716
rect 9124 14682 9158 14716
rect 9192 14682 9226 14716
rect 9260 14682 9294 14716
rect 9328 14682 9362 14716
rect 9396 14682 9430 14716
rect 9464 14682 9498 14716
rect 9532 14682 9566 14716
rect 9674 14688 9708 14722
rect 9742 14688 9776 14722
rect 9810 14688 9844 14722
rect 9926 14682 9960 14716
rect 8964 14566 8998 14600
rect 10050 14606 10084 14640
rect 8964 14498 8998 14532
rect 8964 14430 8998 14464
rect 8964 14362 8998 14396
rect 8964 14294 8998 14328
rect 8964 14226 8998 14260
rect 8964 14158 8998 14192
rect 8964 14090 8998 14124
rect 8964 14022 8998 14056
rect 8964 13954 8998 13988
rect 8964 13886 8998 13920
rect 8964 13818 8998 13852
rect 8964 13750 8998 13784
rect 8964 13682 8998 13716
rect 8964 13614 8998 13648
rect 8890 13522 8924 13556
rect 8964 13546 8998 13580
rect 10050 14538 10084 14572
rect 10050 14470 10084 14504
rect 11470 14628 11504 14662
rect 11538 14628 11572 14662
rect 11606 14628 11640 14662
rect 11674 14628 11708 14662
rect 11742 14628 11776 14662
rect 11810 14628 11844 14662
rect 11878 14628 11912 14662
rect 11946 14628 11980 14662
rect 12014 14628 12048 14662
rect 12082 14628 12116 14662
rect 12150 14628 12184 14662
rect 12218 14628 12252 14662
rect 12286 14628 12320 14662
rect 12354 14628 12388 14662
rect 12422 14628 12456 14662
rect 12490 14628 12524 14662
rect 12558 14628 12592 14662
rect 12626 14628 12660 14662
rect 12694 14628 12728 14662
rect 12762 14628 12796 14662
rect 12830 14628 12864 14662
rect 12898 14628 12932 14662
rect 12966 14628 13000 14662
rect 13034 14628 13068 14662
rect 13102 14628 13136 14662
rect 13170 14628 13204 14662
rect 11446 14517 11480 14551
rect 10050 14402 10084 14436
rect 10050 14334 10084 14368
rect 11446 14449 11480 14483
rect 11446 14381 11480 14415
rect 10050 14266 10084 14300
rect 11446 14313 11480 14347
rect 10050 14198 10084 14232
rect 10050 14130 10084 14164
rect 10050 14062 10084 14096
rect 10050 13994 10084 14028
rect 10050 13926 10084 13960
rect 10050 13858 10084 13892
rect 10050 13790 10084 13824
rect 10050 13722 10084 13756
rect 10050 13654 10084 13688
rect 10050 13553 10084 13587
rect 8866 13417 8900 13451
rect 8866 13349 8900 13383
rect 8866 13281 8900 13315
rect 8866 13213 8900 13247
rect 10050 13485 10084 13519
rect 10050 13417 10084 13451
rect 10050 13349 10084 13383
rect 10050 13281 10084 13315
rect 8940 13189 8974 13223
rect 9008 13189 9042 13223
rect 9076 13189 9110 13223
rect 9144 13189 9178 13223
rect 9212 13189 9246 13223
rect 9280 13189 9314 13223
rect 9348 13189 9382 13223
rect 9372 13058 9406 13092
rect 9372 12990 9406 13024
rect 9372 12922 9406 12956
rect 9372 12854 9406 12888
rect 9372 12786 9406 12820
rect 9372 12718 9406 12752
rect 9372 12650 9406 12684
rect 9372 12582 9406 12616
rect 10050 13213 10084 13247
rect 10050 13145 10084 13179
rect 10050 13077 10084 13111
rect 10050 13009 10084 13043
rect 10050 12941 10084 12975
rect 10050 12873 10084 12907
rect 10050 12805 10084 12839
rect 10050 12737 10084 12771
rect 10050 12669 10084 12703
rect 11446 14245 11480 14279
rect 11446 14177 11480 14211
rect 11446 14109 11480 14143
rect 11446 14041 11480 14075
rect 11446 13973 11480 14007
rect 11446 13905 11480 13939
rect 11446 13837 11480 13871
rect 11446 13769 11480 13803
rect 11446 13701 11480 13735
rect 11446 13633 11480 13667
rect 11446 13565 11480 13599
rect 11446 13497 11480 13531
rect 11446 13429 11480 13463
rect 11446 13361 11480 13395
rect 11446 13293 11480 13327
rect 11446 13225 11480 13259
rect 11446 13157 11480 13191
rect 11446 13089 11480 13123
rect 11446 13021 11480 13055
rect 11446 12953 11480 12987
rect 11446 12885 11480 12919
rect 11446 12784 11480 12818
rect 11446 12716 11480 12750
rect 11446 12648 11480 12682
rect 9343 12433 9377 12467
rect 9343 12365 9377 12399
rect 9343 12297 9377 12331
rect 10079 12534 10113 12568
rect 10079 12466 10113 12500
rect 10079 12398 10113 12432
rect 9443 12273 9477 12307
rect 9511 12273 9545 12307
rect 9579 12273 9613 12307
rect 9647 12273 9681 12307
rect 9715 12273 9749 12307
rect 9783 12273 9817 12307
rect 9851 12273 9885 12307
rect 9919 12273 9953 12307
rect 9987 12273 10021 12307
rect 10055 12273 10089 12307
rect 11446 12580 11480 12614
rect 11446 12512 11480 12546
rect 11446 12444 11480 12478
rect 11446 12376 11480 12410
rect 11446 12308 11480 12342
rect 11446 12240 11480 12274
rect 11446 12172 11480 12206
rect 11446 12104 11480 12138
rect 11446 12036 11480 12070
rect 11446 11968 11480 12002
rect 11446 11900 11480 11934
rect 11446 11832 11480 11866
rect 11446 11764 11480 11798
rect 11446 11696 11480 11730
rect 11446 11628 11480 11662
rect 11446 11560 11480 11594
rect 11446 11492 11480 11526
rect 11446 11424 11480 11458
rect 11446 11356 11480 11390
rect 11446 11288 11480 11322
rect 11446 11220 11480 11254
rect 11446 11152 11480 11186
rect 11446 11084 11480 11118
rect 13254 14604 13288 14638
rect 13254 14536 13288 14570
rect 13254 14468 13288 14502
rect 13254 14400 13288 14434
rect 13254 14332 13288 14366
rect 13254 14264 13288 14298
rect 13254 14196 13288 14230
rect 13254 14128 13288 14162
rect 13254 14060 13288 14094
rect 13254 13992 13288 14026
rect 13254 13924 13288 13958
rect 13254 13856 13288 13890
rect 13254 13788 13288 13822
rect 13254 13720 13288 13754
rect 13254 13652 13288 13686
rect 13254 13584 13288 13618
rect 13254 13516 13288 13550
rect 13254 13448 13288 13482
rect 13254 13380 13288 13414
rect 13254 13312 13288 13346
rect 13254 13244 13288 13278
rect 13254 13176 13288 13210
rect 13342 14604 13376 14638
rect 13434 14628 13468 14662
rect 13502 14628 13536 14662
rect 13570 14628 13604 14662
rect 13638 14628 13672 14662
rect 13706 14628 13740 14662
rect 13774 14628 13808 14662
rect 13842 14628 13876 14662
rect 13910 14628 13944 14662
rect 13978 14628 14012 14662
rect 14046 14628 14080 14662
rect 14114 14628 14148 14662
rect 14182 14628 14216 14662
rect 14250 14628 14284 14662
rect 14318 14628 14352 14662
rect 14386 14628 14420 14662
rect 14454 14628 14488 14662
rect 14522 14628 14556 14662
rect 14590 14628 14624 14662
rect 14658 14628 14692 14662
rect 14726 14628 14760 14662
rect 14794 14628 14828 14662
rect 14862 14628 14896 14662
rect 14930 14628 14964 14662
rect 14998 14628 15032 14662
rect 15066 14628 15100 14662
rect 15134 14628 15168 14662
rect 15202 14628 15236 14662
rect 15270 14628 15304 14662
rect 15338 14628 15372 14662
rect 15406 14628 15440 14662
rect 15474 14628 15508 14662
rect 15542 14628 15576 14662
rect 15610 14628 15644 14662
rect 15678 14628 15712 14662
rect 15746 14628 15780 14662
rect 15814 14628 15848 14662
rect 15882 14628 15916 14662
rect 15950 14628 15984 14662
rect 16018 14628 16052 14662
rect 16086 14628 16120 14662
rect 16154 14628 16188 14662
rect 16222 14628 16256 14662
rect 16290 14628 16324 14662
rect 16358 14628 16392 14662
rect 16426 14628 16460 14662
rect 16494 14628 16528 14662
rect 16562 14628 16596 14662
rect 16630 14628 16664 14662
rect 16698 14628 16732 14662
rect 16766 14628 16800 14662
rect 16834 14628 16868 14662
rect 16902 14628 16936 14662
rect 16970 14628 17004 14662
rect 17038 14628 17072 14662
rect 17106 14628 17140 14662
rect 17174 14628 17208 14662
rect 17242 14628 17276 14662
rect 17310 14628 17344 14662
rect 17378 14628 17412 14662
rect 17446 14628 17480 14662
rect 17514 14628 17548 14662
rect 17582 14628 17616 14662
rect 17650 14628 17684 14662
rect 17718 14628 17752 14662
rect 17786 14628 17820 14662
rect 17854 14628 17888 14662
rect 17922 14628 17956 14662
rect 17990 14628 18024 14662
rect 18058 14628 18092 14662
rect 18126 14628 18160 14662
rect 18194 14628 18228 14662
rect 18262 14628 18296 14662
rect 18330 14628 18364 14662
rect 13342 14536 13376 14570
rect 13342 14468 13376 14502
rect 13342 14400 13376 14434
rect 13342 14332 13376 14366
rect 13342 14264 13376 14298
rect 13342 14196 13376 14230
rect 13342 14128 13376 14162
rect 13342 14060 13376 14094
rect 13342 13992 13376 14026
rect 13342 13924 13376 13958
rect 13342 13856 13376 13890
rect 13342 13788 13376 13822
rect 13342 13720 13376 13754
rect 13342 13652 13376 13686
rect 13342 13584 13376 13618
rect 13342 13516 13376 13550
rect 13342 13448 13376 13482
rect 13342 13380 13376 13414
rect 13342 13312 13376 13346
rect 13342 13244 13376 13278
rect 18354 14560 18388 14594
rect 18354 14492 18388 14526
rect 18354 14424 18388 14458
rect 18354 14356 18388 14390
rect 18354 14288 18388 14322
rect 18354 14220 18388 14254
rect 18354 14152 18388 14186
rect 18354 14084 18388 14118
rect 18354 14016 18388 14050
rect 18354 13948 18388 13982
rect 18354 13880 18388 13914
rect 18354 13812 18388 13846
rect 18354 13744 18388 13778
rect 18354 13676 18388 13710
rect 18354 13608 18388 13642
rect 18354 13540 18388 13574
rect 18354 13472 18388 13506
rect 18354 13404 18388 13438
rect 18354 13336 18388 13370
rect 18354 13268 18388 13302
rect 13366 13176 13400 13210
rect 13434 13176 13468 13210
rect 13502 13176 13536 13210
rect 13570 13176 13604 13210
rect 13638 13176 13672 13210
rect 13706 13176 13740 13210
rect 13774 13176 13808 13210
rect 13842 13176 13876 13210
rect 13910 13176 13944 13210
rect 13978 13176 14012 13210
rect 14046 13176 14080 13210
rect 14114 13176 14148 13210
rect 14182 13176 14216 13210
rect 14250 13176 14284 13210
rect 14318 13176 14352 13210
rect 14386 13176 14420 13210
rect 14454 13176 14488 13210
rect 14522 13176 14556 13210
rect 14590 13176 14624 13210
rect 14658 13176 14692 13210
rect 14726 13176 14760 13210
rect 14794 13176 14828 13210
rect 14862 13176 14896 13210
rect 14930 13176 14964 13210
rect 14998 13176 15032 13210
rect 15066 13176 15100 13210
rect 15134 13176 15168 13210
rect 15202 13176 15236 13210
rect 15270 13176 15304 13210
rect 15338 13176 15372 13210
rect 15406 13176 15440 13210
rect 15474 13176 15508 13210
rect 15542 13176 15576 13210
rect 15610 13176 15644 13210
rect 15678 13176 15712 13210
rect 15746 13176 15780 13210
rect 15889 13176 15923 13210
rect 15957 13176 15991 13210
rect 16025 13176 16059 13210
rect 16093 13176 16127 13210
rect 16161 13176 16195 13210
rect 16229 13176 16263 13210
rect 16297 13176 16331 13210
rect 16365 13176 16399 13210
rect 16433 13176 16467 13210
rect 16501 13176 16535 13210
rect 16569 13176 16603 13210
rect 16637 13176 16671 13210
rect 16705 13176 16739 13210
rect 16773 13176 16807 13210
rect 16841 13176 16875 13210
rect 16909 13176 16943 13210
rect 16977 13176 17011 13210
rect 17045 13176 17079 13210
rect 17113 13176 17147 13210
rect 17181 13176 17215 13210
rect 17249 13176 17283 13210
rect 17317 13176 17351 13210
rect 17385 13176 17419 13210
rect 17453 13176 17487 13210
rect 17521 13176 17555 13210
rect 17589 13176 17623 13210
rect 17657 13176 17691 13210
rect 17725 13176 17759 13210
rect 17793 13176 17827 13210
rect 17861 13176 17895 13210
rect 17929 13176 17963 13210
rect 17997 13176 18031 13210
rect 18065 13176 18099 13210
rect 18133 13176 18167 13210
rect 18201 13176 18235 13210
rect 18269 13176 18303 13210
rect 18354 13200 18388 13234
rect 13254 13108 13288 13142
rect 13254 13040 13288 13074
rect 13254 12972 13288 13006
rect 13254 12904 13288 12938
rect 13254 12836 13288 12870
rect 13254 12768 13288 12802
rect 13254 12700 13288 12734
rect 13254 12632 13288 12666
rect 13254 12564 13288 12598
rect 13254 12496 13288 12530
rect 13254 12428 13288 12462
rect 13254 12360 13288 12394
rect 13254 12292 13288 12326
rect 13254 12224 13288 12258
rect 13254 12156 13288 12190
rect 13254 12088 13288 12122
rect 13254 12020 13288 12054
rect 13254 11952 13288 11986
rect 13254 11884 13288 11918
rect 13254 11816 13288 11850
rect 13254 11748 13288 11782
rect 13254 11680 13288 11714
rect 13254 11612 13288 11646
rect 13254 11544 13288 11578
rect 13254 11476 13288 11510
rect 13254 11408 13288 11442
rect 13254 11340 13288 11374
rect 13254 11272 13288 11306
rect 13254 11204 13288 11238
rect 13254 11136 13288 11170
rect 11530 11060 11564 11094
rect 11598 11060 11632 11094
rect 11666 11060 11700 11094
rect 11734 11060 11768 11094
rect 11802 11060 11836 11094
rect 11870 11060 11904 11094
rect 11938 11060 11972 11094
rect 12006 11060 12040 11094
rect 12074 11060 12108 11094
rect 12142 11060 12176 11094
rect 12210 11060 12244 11094
rect 12278 11060 12312 11094
rect 12346 11060 12380 11094
rect 12414 11060 12448 11094
rect 12482 11060 12516 11094
rect 12550 11060 12584 11094
rect 12618 11060 12652 11094
rect 12686 11060 12720 11094
rect 12754 11060 12788 11094
rect 12822 11060 12856 11094
rect 12890 11060 12924 11094
rect 12958 11060 12992 11094
rect 13026 11060 13060 11094
rect 13094 11060 13128 11094
rect 13162 11060 13196 11094
rect 13230 11060 13264 11094
<< nsubdiffcont >>
rect 9469 37602 9503 37636
rect 9537 37602 9571 37636
rect 9605 37602 9639 37636
rect 9673 37602 9707 37636
rect 9741 37602 9775 37636
rect 9809 37602 9843 37636
rect 9877 37602 9911 37636
rect 9945 37602 9979 37636
rect 10013 37602 10047 37636
rect 10081 37602 10115 37636
rect 10149 37602 10183 37636
rect 10217 37602 10251 37636
rect 10285 37602 10319 37636
rect 10353 37602 10387 37636
rect 10421 37602 10455 37636
rect 10489 37602 10523 37636
rect 10557 37602 10591 37636
rect 10625 37602 10659 37636
rect 10693 37602 10727 37636
rect 10761 37602 10795 37636
rect 10829 37602 10863 37636
rect 10897 37602 10931 37636
rect 10965 37602 10999 37636
rect 11033 37602 11067 37636
rect 11101 37602 11135 37636
rect 11169 37602 11203 37636
rect 11237 37602 11271 37636
rect 11305 37602 11339 37636
rect 11373 37602 11407 37636
rect 11441 37602 11475 37636
rect 11509 37602 11543 37636
rect 11577 37602 11611 37636
rect 11645 37602 11679 37636
rect 11713 37602 11747 37636
rect 11781 37602 11815 37636
rect 11849 37602 11883 37636
rect 11917 37602 11951 37636
rect 11985 37602 12019 37636
rect 12053 37602 12087 37636
rect 12121 37602 12155 37636
rect 12189 37602 12223 37636
rect 12257 37602 12291 37636
rect 12348 37602 12382 37636
rect 12416 37602 12450 37636
rect 12484 37602 12518 37636
rect 12552 37602 12586 37636
rect 12620 37602 12654 37636
rect 12688 37602 12722 37636
rect 12756 37602 12790 37636
rect 12824 37602 12858 37636
rect 12892 37602 12926 37636
rect 12960 37602 12994 37636
rect 13028 37602 13062 37636
rect 13096 37602 13130 37636
rect 13164 37602 13198 37636
rect 13232 37602 13266 37636
rect 13300 37602 13334 37636
rect 13368 37602 13402 37636
rect 13436 37602 13470 37636
rect 13504 37602 13538 37636
rect 13572 37602 13606 37636
rect 13640 37602 13674 37636
rect 13708 37602 13742 37636
rect 13776 37602 13810 37636
rect 13844 37602 13878 37636
rect 13912 37602 13946 37636
rect 13980 37602 14014 37636
rect 14048 37602 14082 37636
rect 14116 37602 14150 37636
rect 14184 37602 14218 37636
rect 14252 37602 14286 37636
rect 14320 37602 14354 37636
rect 14388 37602 14422 37636
rect 14456 37602 14490 37636
rect 14524 37602 14558 37636
rect 14592 37602 14626 37636
rect 14660 37602 14694 37636
rect 14728 37602 14762 37636
rect 14796 37602 14830 37636
rect 14864 37602 14898 37636
rect 14932 37602 14966 37636
rect 15000 37602 15034 37636
rect 15068 37602 15102 37636
rect 9445 37508 9479 37542
rect 15169 37578 15203 37612
rect 9445 37440 9479 37474
rect 9599 37466 9633 37500
rect 9667 37466 9701 37500
rect 9735 37466 9769 37500
rect 9803 37466 9837 37500
rect 9871 37466 9905 37500
rect 9939 37466 9973 37500
rect 10007 37466 10041 37500
rect 10075 37466 10109 37500
rect 10143 37466 10177 37500
rect 10211 37466 10245 37500
rect 10374 37466 10408 37500
rect 10442 37466 10476 37500
rect 10510 37466 10544 37500
rect 10578 37466 10612 37500
rect 10646 37466 10680 37500
rect 10714 37466 10748 37500
rect 10782 37466 10816 37500
rect 10850 37466 10884 37500
rect 10918 37466 10952 37500
rect 11034 37466 11068 37500
rect 11102 37466 11136 37500
rect 11170 37466 11204 37500
rect 11238 37466 11272 37500
rect 11306 37466 11340 37500
rect 11374 37466 11408 37500
rect 11442 37466 11476 37500
rect 11510 37466 11544 37500
rect 11578 37466 11612 37500
rect 11690 37466 11724 37500
rect 11758 37466 11792 37500
rect 11826 37466 11860 37500
rect 11894 37466 11928 37500
rect 11962 37466 11996 37500
rect 12030 37466 12064 37500
rect 12098 37466 12132 37500
rect 12166 37466 12200 37500
rect 12234 37466 12268 37500
rect 12363 37466 12397 37500
rect 12431 37466 12465 37500
rect 12499 37466 12533 37500
rect 12567 37466 12601 37500
rect 12635 37466 12669 37500
rect 12703 37466 12737 37500
rect 12771 37466 12805 37500
rect 12839 37466 12873 37500
rect 12907 37466 12941 37500
rect 13036 37466 13070 37500
rect 13104 37466 13138 37500
rect 13172 37466 13206 37500
rect 13240 37466 13274 37500
rect 13308 37466 13342 37500
rect 13376 37466 13410 37500
rect 13444 37466 13478 37500
rect 13512 37466 13546 37500
rect 13580 37466 13614 37500
rect 13696 37466 13730 37500
rect 13764 37466 13798 37500
rect 13832 37466 13866 37500
rect 13900 37466 13934 37500
rect 13968 37466 14002 37500
rect 14036 37466 14070 37500
rect 14104 37466 14138 37500
rect 14172 37466 14206 37500
rect 14240 37466 14274 37500
rect 15169 37510 15203 37544
rect 15169 37442 15203 37476
rect 9445 37372 9479 37406
rect 9445 37304 9479 37338
rect 9445 37236 9479 37270
rect 9445 37168 9479 37202
rect 9445 37100 9479 37134
rect 9445 37032 9479 37066
rect 9445 36964 9479 36998
rect 9445 36896 9479 36930
rect 9445 36828 9479 36862
rect 9445 36760 9479 36794
rect 9445 36692 9479 36726
rect 9445 36624 9479 36658
rect 9445 36556 9479 36590
rect 9445 36488 9479 36522
rect 9445 36420 9479 36454
rect 9445 36352 9479 36386
rect 9445 36284 9479 36318
rect 9445 36216 9479 36250
rect 9445 36148 9479 36182
rect 9445 36080 9479 36114
rect 9445 36012 9479 36046
rect 15169 37374 15203 37408
rect 15169 37306 15203 37340
rect 15169 37238 15203 37272
rect 15169 37170 15203 37204
rect 15169 37102 15203 37136
rect 15169 37034 15203 37068
rect 15169 36966 15203 37000
rect 15169 36898 15203 36932
rect 15169 36830 15203 36864
rect 15169 36762 15203 36796
rect 15169 36694 15203 36728
rect 15169 36626 15203 36660
rect 15169 36558 15203 36592
rect 15169 36490 15203 36524
rect 15169 36422 15203 36456
rect 15169 36354 15203 36388
rect 15169 36286 15203 36320
rect 15169 36218 15203 36252
rect 15169 36150 15203 36184
rect 15169 36082 15203 36116
rect 9445 35944 9479 35978
rect 15169 36014 15203 36048
rect 9445 35876 9479 35910
rect 9445 35808 9479 35842
rect 9445 35740 9479 35774
rect 9445 35672 9479 35706
rect 9445 35604 9479 35638
rect 9445 35536 9479 35570
rect 9445 35468 9479 35502
rect 9445 35400 9479 35434
rect 9445 35332 9479 35366
rect 9445 35264 9479 35298
rect 9445 35196 9479 35230
rect 9445 35128 9479 35162
rect 9445 35060 9479 35094
rect 9445 34992 9479 35026
rect 9445 34924 9479 34958
rect 9445 34856 9479 34890
rect 9445 34788 9479 34822
rect 6976 34688 7010 34722
rect 7044 34688 7078 34722
rect 7112 34688 7146 34722
rect 7180 34688 7214 34722
rect 7248 34688 7282 34722
rect 7316 34688 7350 34722
rect 7384 34688 7418 34722
rect 7452 34688 7486 34722
rect 7520 34688 7554 34722
rect 7588 34688 7622 34722
rect 7656 34688 7690 34722
rect 7724 34688 7758 34722
rect 7792 34688 7826 34722
rect 6952 34608 6986 34642
rect 6952 34540 6986 34574
rect 6952 34472 6986 34506
rect 6952 34404 6986 34438
rect 6952 34336 6986 34370
rect 6952 34268 6986 34302
rect 6952 34200 6986 34234
rect 6952 34132 6986 34166
rect 6952 34064 6986 34098
rect 6952 33996 6986 34030
rect 6952 33857 6986 33891
rect 6952 33789 6986 33823
rect 6952 33721 6986 33755
rect 6952 33653 6986 33687
rect 6952 33585 6986 33619
rect 6952 33517 6986 33551
rect 6952 33449 6986 33483
rect 6952 33381 6986 33415
rect 6952 33313 6986 33347
rect 6952 33245 6986 33279
rect 7892 34664 7926 34698
rect 7892 34596 7926 34630
rect 7892 34528 7926 34562
rect 7892 34460 7926 34494
rect 7892 34392 7926 34426
rect 9445 34720 9479 34754
rect 9445 34652 9479 34686
rect 9445 34584 9479 34618
rect 15169 35946 15203 35980
rect 15169 35878 15203 35912
rect 15169 35810 15203 35844
rect 15169 35742 15203 35776
rect 15169 35674 15203 35708
rect 15169 35606 15203 35640
rect 15169 35538 15203 35572
rect 15169 35470 15203 35504
rect 15169 35402 15203 35436
rect 15169 35334 15203 35368
rect 15169 35266 15203 35300
rect 15169 35198 15203 35232
rect 15169 35130 15203 35164
rect 15169 35062 15203 35096
rect 15169 34994 15203 35028
rect 15169 34926 15203 34960
rect 15169 34858 15203 34892
rect 15169 34790 15203 34824
rect 15169 34722 15203 34756
rect 15169 34654 15203 34688
rect 9445 34516 9479 34550
rect 15169 34586 15203 34620
rect 9445 34448 9479 34482
rect 15169 34518 15203 34552
rect 9569 34424 9603 34458
rect 9637 34424 9671 34458
rect 9705 34424 9739 34458
rect 9773 34424 9807 34458
rect 9841 34424 9875 34458
rect 9909 34424 9943 34458
rect 9977 34424 10011 34458
rect 10045 34424 10079 34458
rect 10113 34424 10147 34458
rect 10181 34424 10215 34458
rect 10249 34424 10283 34458
rect 10317 34424 10351 34458
rect 10385 34424 10419 34458
rect 10453 34424 10487 34458
rect 10521 34424 10555 34458
rect 10589 34424 10623 34458
rect 10657 34424 10691 34458
rect 10725 34424 10759 34458
rect 10793 34424 10827 34458
rect 10861 34424 10895 34458
rect 10929 34424 10963 34458
rect 10997 34424 11031 34458
rect 11065 34424 11099 34458
rect 11133 34424 11167 34458
rect 11201 34424 11235 34458
rect 11269 34424 11303 34458
rect 11337 34424 11371 34458
rect 11405 34424 11439 34458
rect 11473 34424 11507 34458
rect 11541 34424 11575 34458
rect 11609 34424 11643 34458
rect 11677 34424 11711 34458
rect 11745 34424 11779 34458
rect 11813 34424 11847 34458
rect 11881 34424 11915 34458
rect 11949 34424 11983 34458
rect 12017 34424 12051 34458
rect 12085 34424 12119 34458
rect 12153 34424 12187 34458
rect 12221 34424 12255 34458
rect 12289 34424 12323 34458
rect 12357 34424 12391 34458
rect 12425 34424 12459 34458
rect 12493 34424 12527 34458
rect 12561 34424 12595 34458
rect 12629 34424 12663 34458
rect 12697 34424 12731 34458
rect 12765 34424 12799 34458
rect 12833 34424 12867 34458
rect 12901 34424 12935 34458
rect 12969 34424 13003 34458
rect 13037 34424 13071 34458
rect 13105 34424 13139 34458
rect 13173 34424 13207 34458
rect 13241 34424 13275 34458
rect 13309 34424 13343 34458
rect 13377 34424 13411 34458
rect 13445 34424 13479 34458
rect 13513 34424 13547 34458
rect 13581 34424 13615 34458
rect 13649 34424 13683 34458
rect 13717 34424 13751 34458
rect 13785 34424 13819 34458
rect 13853 34424 13887 34458
rect 13921 34424 13955 34458
rect 13989 34424 14023 34458
rect 14057 34424 14091 34458
rect 14125 34424 14159 34458
rect 14193 34424 14227 34458
rect 14261 34424 14295 34458
rect 14329 34424 14363 34458
rect 14397 34424 14431 34458
rect 14465 34424 14499 34458
rect 14533 34424 14567 34458
rect 14601 34424 14635 34458
rect 14669 34424 14703 34458
rect 14737 34424 14771 34458
rect 14805 34424 14839 34458
rect 14873 34424 14907 34458
rect 14941 34424 14975 34458
rect 15009 34424 15043 34458
rect 15077 34424 15111 34458
rect 15145 34424 15179 34458
rect 15275 37578 15309 37612
rect 15371 37602 15405 37636
rect 15439 37602 15473 37636
rect 15507 37602 15541 37636
rect 15575 37602 15609 37636
rect 15643 37602 15677 37636
rect 15711 37602 15745 37636
rect 15779 37602 15813 37636
rect 15847 37602 15881 37636
rect 15915 37602 15949 37636
rect 15983 37602 16017 37636
rect 16051 37602 16085 37636
rect 16119 37602 16153 37636
rect 16187 37602 16221 37636
rect 16255 37602 16289 37636
rect 16323 37602 16357 37636
rect 16391 37602 16425 37636
rect 16459 37602 16493 37636
rect 16527 37602 16561 37636
rect 16595 37602 16629 37636
rect 16663 37602 16697 37636
rect 16731 37602 16765 37636
rect 16799 37602 16833 37636
rect 16867 37602 16901 37636
rect 16935 37602 16969 37636
rect 17003 37602 17037 37636
rect 17071 37602 17105 37636
rect 17139 37602 17173 37636
rect 17207 37602 17241 37636
rect 17275 37602 17309 37636
rect 17343 37602 17377 37636
rect 17411 37602 17445 37636
rect 17479 37602 17513 37636
rect 17547 37602 17581 37636
rect 17615 37602 17649 37636
rect 17683 37602 17717 37636
rect 17751 37602 17785 37636
rect 17819 37602 17853 37636
rect 17887 37602 17921 37636
rect 17955 37602 17989 37636
rect 18023 37602 18057 37636
rect 18091 37602 18125 37636
rect 18159 37602 18193 37636
rect 15275 37510 15309 37544
rect 15275 37442 15309 37476
rect 15275 37374 15309 37408
rect 15275 37306 15309 37340
rect 15275 37238 15309 37272
rect 15275 37170 15309 37204
rect 15275 37102 15309 37136
rect 15275 37034 15309 37068
rect 15275 36966 15309 37000
rect 15275 36898 15309 36932
rect 15275 36830 15309 36864
rect 15275 36762 15309 36796
rect 15275 36694 15309 36728
rect 15275 36626 15309 36660
rect 15275 36558 15309 36592
rect 15275 36490 15309 36524
rect 15275 36422 15309 36456
rect 15275 36354 15309 36388
rect 15275 36286 15309 36320
rect 15275 36218 15309 36252
rect 15275 36150 15309 36184
rect 15275 36082 15309 36116
rect 15275 36014 15309 36048
rect 15275 35946 15309 35980
rect 15275 35878 15309 35912
rect 15275 35810 15309 35844
rect 15275 35742 15309 35776
rect 15275 35674 15309 35708
rect 15275 35606 15309 35640
rect 15275 35538 15309 35572
rect 15275 35470 15309 35504
rect 15275 35402 15309 35436
rect 15275 35334 15309 35368
rect 15275 35266 15309 35300
rect 15275 35198 15309 35232
rect 15275 35130 15309 35164
rect 15275 35062 15309 35096
rect 15275 34994 15309 35028
rect 15275 34926 15309 34960
rect 15275 34858 15309 34892
rect 15275 34790 15309 34824
rect 15275 34722 15309 34756
rect 15275 34654 15309 34688
rect 15275 34586 15309 34620
rect 15275 34518 15309 34552
rect 18183 37482 18217 37516
rect 18183 37414 18217 37448
rect 18183 37346 18217 37380
rect 18183 37278 18217 37312
rect 18183 37210 18217 37244
rect 18183 37142 18217 37176
rect 18183 37074 18217 37108
rect 18183 37006 18217 37040
rect 18183 36938 18217 36972
rect 18183 36870 18217 36904
rect 18183 36802 18217 36836
rect 18183 36734 18217 36768
rect 18183 36666 18217 36700
rect 18183 36598 18217 36632
rect 18183 36530 18217 36564
rect 18183 36462 18217 36496
rect 18183 36394 18217 36428
rect 18183 36326 18217 36360
rect 18183 36258 18217 36292
rect 18183 36190 18217 36224
rect 18183 36122 18217 36156
rect 18183 36054 18217 36088
rect 18183 35944 18217 35978
rect 18183 35876 18217 35910
rect 18183 35808 18217 35842
rect 18183 35740 18217 35774
rect 18183 35672 18217 35706
rect 18183 35604 18217 35638
rect 18183 35536 18217 35570
rect 18183 35468 18217 35502
rect 18183 35400 18217 35434
rect 18183 35332 18217 35366
rect 18183 35264 18217 35298
rect 18183 35196 18217 35230
rect 18183 35128 18217 35162
rect 18183 35060 18217 35094
rect 18183 34992 18217 35026
rect 18183 34924 18217 34958
rect 18183 34856 18217 34890
rect 18183 34788 18217 34822
rect 18183 34720 18217 34754
rect 18183 34652 18217 34686
rect 18183 34584 18217 34618
rect 18183 34516 18217 34550
rect 15299 34424 15333 34458
rect 15367 34424 15401 34458
rect 15435 34424 15469 34458
rect 15503 34424 15537 34458
rect 15571 34424 15605 34458
rect 15639 34424 15673 34458
rect 15707 34424 15741 34458
rect 15775 34424 15809 34458
rect 15843 34424 15877 34458
rect 15911 34424 15945 34458
rect 15979 34424 16013 34458
rect 16047 34424 16081 34458
rect 16115 34424 16149 34458
rect 16183 34424 16217 34458
rect 16251 34424 16285 34458
rect 16319 34424 16353 34458
rect 16387 34424 16421 34458
rect 16455 34424 16489 34458
rect 16523 34424 16557 34458
rect 16591 34424 16625 34458
rect 16659 34424 16693 34458
rect 16727 34424 16761 34458
rect 16795 34424 16829 34458
rect 16863 34424 16897 34458
rect 16931 34424 16965 34458
rect 16999 34424 17033 34458
rect 17067 34424 17101 34458
rect 17135 34424 17169 34458
rect 17203 34424 17237 34458
rect 17271 34424 17305 34458
rect 17339 34424 17373 34458
rect 17407 34424 17441 34458
rect 17475 34424 17509 34458
rect 17543 34424 17577 34458
rect 17611 34424 17645 34458
rect 17679 34424 17713 34458
rect 17747 34424 17781 34458
rect 17815 34424 17849 34458
rect 17883 34424 17917 34458
rect 17951 34424 17985 34458
rect 18019 34424 18053 34458
rect 18087 34424 18121 34458
rect 18183 34448 18217 34482
rect 18289 37578 18323 37612
rect 18362 37602 18396 37636
rect 18430 37602 18464 37636
rect 18498 37602 18532 37636
rect 18566 37602 18600 37636
rect 18634 37602 18668 37636
rect 18702 37602 18736 37636
rect 18770 37602 18804 37636
rect 18838 37602 18872 37636
rect 18906 37602 18940 37636
rect 18974 37602 19008 37636
rect 19042 37602 19076 37636
rect 19110 37602 19144 37636
rect 19178 37602 19212 37636
rect 19246 37602 19280 37636
rect 19314 37602 19348 37636
rect 19382 37602 19416 37636
rect 19450 37602 19484 37636
rect 19518 37602 19552 37636
rect 19586 37602 19620 37636
rect 19654 37602 19688 37636
rect 19722 37602 19756 37636
rect 19790 37602 19824 37636
rect 19858 37602 19892 37636
rect 19926 37602 19960 37636
rect 19994 37602 20028 37636
rect 20062 37602 20096 37636
rect 20130 37602 20164 37636
rect 20198 37602 20232 37636
rect 20266 37602 20300 37636
rect 20334 37602 20368 37636
rect 20402 37602 20436 37636
rect 20470 37602 20504 37636
rect 20538 37602 20572 37636
rect 20606 37602 20640 37636
rect 20674 37602 20708 37636
rect 20742 37602 20776 37636
rect 20810 37602 20844 37636
rect 20878 37602 20912 37636
rect 20946 37602 20980 37636
rect 21014 37602 21048 37636
rect 21145 37602 21179 37636
rect 21213 37602 21247 37636
rect 21281 37602 21315 37636
rect 21349 37602 21383 37636
rect 21417 37602 21451 37636
rect 21485 37602 21519 37636
rect 21553 37602 21587 37636
rect 21621 37602 21655 37636
rect 21689 37602 21723 37636
rect 21757 37602 21791 37636
rect 21825 37602 21859 37636
rect 21893 37602 21927 37636
rect 21961 37602 21995 37636
rect 22029 37602 22063 37636
rect 22097 37602 22131 37636
rect 22165 37602 22199 37636
rect 22233 37602 22267 37636
rect 22301 37602 22335 37636
rect 22369 37602 22403 37636
rect 22437 37602 22471 37636
rect 22505 37602 22539 37636
rect 22573 37602 22607 37636
rect 22641 37602 22675 37636
rect 22709 37602 22743 37636
rect 22777 37602 22811 37636
rect 22845 37602 22879 37636
rect 22913 37602 22947 37636
rect 22981 37602 23015 37636
rect 23049 37602 23083 37636
rect 23117 37602 23151 37636
rect 23185 37602 23219 37636
rect 23253 37602 23287 37636
rect 23321 37602 23355 37636
rect 23389 37602 23423 37636
rect 23457 37602 23491 37636
rect 23525 37602 23559 37636
rect 23593 37602 23627 37636
rect 23661 37602 23695 37636
rect 23729 37602 23763 37636
rect 23797 37602 23831 37636
rect 18289 37510 18323 37544
rect 23821 37508 23855 37542
rect 18289 37442 18323 37476
rect 19143 37448 19177 37482
rect 19211 37448 19245 37482
rect 19279 37448 19313 37482
rect 19347 37448 19381 37482
rect 19415 37448 19449 37482
rect 19483 37448 19517 37482
rect 19551 37448 19585 37482
rect 19619 37448 19653 37482
rect 19687 37448 19721 37482
rect 19816 37448 19850 37482
rect 19884 37448 19918 37482
rect 19952 37448 19986 37482
rect 20020 37448 20054 37482
rect 20088 37448 20122 37482
rect 20156 37448 20190 37482
rect 20224 37448 20258 37482
rect 20292 37448 20326 37482
rect 20360 37448 20394 37482
rect 20489 37448 20523 37482
rect 20557 37448 20591 37482
rect 20625 37448 20659 37482
rect 20693 37448 20727 37482
rect 20761 37448 20795 37482
rect 20829 37448 20863 37482
rect 20897 37448 20931 37482
rect 20965 37448 20999 37482
rect 21094 37448 21128 37482
rect 21162 37448 21196 37482
rect 21230 37448 21264 37482
rect 21298 37448 21332 37482
rect 21366 37448 21400 37482
rect 21434 37448 21468 37482
rect 21502 37448 21536 37482
rect 21570 37448 21604 37482
rect 21638 37448 21672 37482
rect 21767 37448 21801 37482
rect 21835 37448 21869 37482
rect 21903 37448 21937 37482
rect 21971 37448 22005 37482
rect 22039 37448 22073 37482
rect 22107 37448 22141 37482
rect 22175 37448 22209 37482
rect 22243 37448 22277 37482
rect 22311 37448 22345 37482
rect 22440 37448 22474 37482
rect 22508 37448 22542 37482
rect 22576 37448 22610 37482
rect 22644 37448 22678 37482
rect 22712 37448 22746 37482
rect 22780 37448 22814 37482
rect 22848 37448 22882 37482
rect 22916 37448 22950 37482
rect 22984 37448 23018 37482
rect 23821 37440 23855 37474
rect 18289 37374 18323 37408
rect 23821 37372 23855 37406
rect 18289 37306 18323 37340
rect 18289 37238 18323 37272
rect 18289 37170 18323 37204
rect 18289 37102 18323 37136
rect 18289 37034 18323 37068
rect 18289 36966 18323 37000
rect 18289 36898 18323 36932
rect 18289 36830 18323 36864
rect 18289 36762 18323 36796
rect 18289 36694 18323 36728
rect 18289 36626 18323 36660
rect 18289 36558 18323 36592
rect 18289 36490 18323 36524
rect 18289 36422 18323 36456
rect 18289 36354 18323 36388
rect 18289 36286 18323 36320
rect 18289 36218 18323 36252
rect 18289 36150 18323 36184
rect 18289 36082 18323 36116
rect 18289 36014 18323 36048
rect 23821 37304 23855 37338
rect 23821 37236 23855 37270
rect 23821 37168 23855 37202
rect 23821 37100 23855 37134
rect 23821 37032 23855 37066
rect 23821 36964 23855 36998
rect 23821 36896 23855 36930
rect 23821 36828 23855 36862
rect 23821 36760 23855 36794
rect 23821 36692 23855 36726
rect 23821 36624 23855 36658
rect 23821 36556 23855 36590
rect 23821 36488 23855 36522
rect 23821 36420 23855 36454
rect 23821 36352 23855 36386
rect 23821 36284 23855 36318
rect 23821 36216 23855 36250
rect 23821 36148 23855 36182
rect 23821 36080 23855 36114
rect 23821 36012 23855 36046
rect 18289 35946 18323 35980
rect 18289 35878 18323 35912
rect 18289 35810 18323 35844
rect 18289 35742 18323 35776
rect 18289 35674 18323 35708
rect 18289 35606 18323 35640
rect 18289 35538 18323 35572
rect 18289 35470 18323 35504
rect 18289 35402 18323 35436
rect 18289 35334 18323 35368
rect 18289 35266 18323 35300
rect 18289 35198 18323 35232
rect 18289 35130 18323 35164
rect 18289 35062 18323 35096
rect 18289 34994 18323 35028
rect 18289 34926 18323 34960
rect 18289 34858 18323 34892
rect 18289 34790 18323 34824
rect 18289 34722 18323 34756
rect 18289 34654 18323 34688
rect 18289 34586 18323 34620
rect 18289 34518 18323 34552
rect 23821 35944 23855 35978
rect 23821 35876 23855 35910
rect 23821 35808 23855 35842
rect 23821 35740 23855 35774
rect 23821 35672 23855 35706
rect 23821 35604 23855 35638
rect 23821 35536 23855 35570
rect 23821 35468 23855 35502
rect 23821 35400 23855 35434
rect 23821 35332 23855 35366
rect 23821 35264 23855 35298
rect 23821 35196 23855 35230
rect 23821 35128 23855 35162
rect 23821 35060 23855 35094
rect 23821 34992 23855 35026
rect 23821 34924 23855 34958
rect 23821 34856 23855 34890
rect 23821 34788 23855 34822
rect 23821 34720 23855 34754
rect 23821 34652 23855 34686
rect 23821 34584 23855 34618
rect 23821 34516 23855 34550
rect 18313 34424 18347 34458
rect 18381 34424 18415 34458
rect 18449 34424 18483 34458
rect 18517 34424 18551 34458
rect 18585 34424 18619 34458
rect 18653 34424 18687 34458
rect 18721 34424 18755 34458
rect 18789 34424 18823 34458
rect 18857 34424 18891 34458
rect 18925 34424 18959 34458
rect 18993 34424 19027 34458
rect 19061 34424 19095 34458
rect 19129 34424 19163 34458
rect 19197 34424 19231 34458
rect 19265 34424 19299 34458
rect 19333 34424 19367 34458
rect 19401 34424 19435 34458
rect 19469 34424 19503 34458
rect 19537 34424 19571 34458
rect 19605 34424 19639 34458
rect 19673 34424 19707 34458
rect 19741 34424 19775 34458
rect 19809 34424 19843 34458
rect 19877 34424 19911 34458
rect 19945 34424 19979 34458
rect 20013 34424 20047 34458
rect 20081 34424 20115 34458
rect 20149 34424 20183 34458
rect 20217 34424 20251 34458
rect 20285 34424 20319 34458
rect 20353 34424 20387 34458
rect 20421 34424 20455 34458
rect 20489 34424 20523 34458
rect 20557 34424 20591 34458
rect 20625 34424 20659 34458
rect 20693 34424 20727 34458
rect 20761 34424 20795 34458
rect 20829 34424 20863 34458
rect 20897 34424 20931 34458
rect 20965 34424 20999 34458
rect 21033 34424 21067 34458
rect 21101 34424 21135 34458
rect 21169 34424 21203 34458
rect 21237 34424 21271 34458
rect 21305 34424 21339 34458
rect 21373 34424 21407 34458
rect 21441 34424 21475 34458
rect 21509 34424 21543 34458
rect 21577 34424 21611 34458
rect 21645 34424 21679 34458
rect 21713 34424 21747 34458
rect 21781 34424 21815 34458
rect 21849 34424 21883 34458
rect 21917 34424 21951 34458
rect 21985 34424 22019 34458
rect 22053 34424 22087 34458
rect 22121 34424 22155 34458
rect 22189 34424 22223 34458
rect 22257 34424 22291 34458
rect 22325 34424 22359 34458
rect 22393 34424 22427 34458
rect 22461 34424 22495 34458
rect 22529 34424 22563 34458
rect 22597 34424 22631 34458
rect 22665 34424 22699 34458
rect 22733 34424 22767 34458
rect 22801 34424 22835 34458
rect 22869 34424 22903 34458
rect 22937 34424 22971 34458
rect 23005 34424 23039 34458
rect 23073 34424 23107 34458
rect 23141 34424 23175 34458
rect 23209 34424 23243 34458
rect 23277 34424 23311 34458
rect 23345 34424 23379 34458
rect 23413 34424 23447 34458
rect 23481 34424 23515 34458
rect 23549 34424 23583 34458
rect 23617 34424 23651 34458
rect 23685 34424 23719 34458
rect 23753 34424 23787 34458
rect 23821 34448 23855 34482
rect 7892 34324 7926 34358
rect 7892 34256 7926 34290
rect 7892 34188 7926 34222
rect 7892 34120 7926 34154
rect 7892 34052 7926 34086
rect 7892 33984 7926 34018
rect 7892 33916 7926 33950
rect 7892 33848 7926 33882
rect 7892 33780 7926 33814
rect 7892 33712 7926 33746
rect 7892 33644 7926 33678
rect 9469 34318 9503 34352
rect 9537 34318 9571 34352
rect 9605 34318 9639 34352
rect 9673 34318 9707 34352
rect 9741 34318 9775 34352
rect 9809 34318 9843 34352
rect 9877 34318 9911 34352
rect 9945 34318 9979 34352
rect 10013 34318 10047 34352
rect 10081 34318 10115 34352
rect 10149 34318 10183 34352
rect 10217 34318 10251 34352
rect 10285 34318 10319 34352
rect 10353 34318 10387 34352
rect 10421 34318 10455 34352
rect 10489 34318 10523 34352
rect 10637 34318 10671 34352
rect 10705 34318 10739 34352
rect 10773 34318 10807 34352
rect 10841 34318 10875 34352
rect 10909 34318 10943 34352
rect 10977 34318 11011 34352
rect 11045 34318 11079 34352
rect 11113 34318 11147 34352
rect 11181 34318 11215 34352
rect 11249 34318 11283 34352
rect 11317 34318 11351 34352
rect 11385 34318 11419 34352
rect 11453 34318 11487 34352
rect 11521 34318 11555 34352
rect 11589 34318 11623 34352
rect 11657 34318 11691 34352
rect 9445 34244 9479 34278
rect 9445 34176 9479 34210
rect 11747 34294 11781 34328
rect 11747 34226 11781 34260
rect 9445 34108 9479 34142
rect 11747 34158 11781 34192
rect 9445 34040 9479 34074
rect 9445 33972 9479 34006
rect 9445 33904 9479 33938
rect 9445 33836 9479 33870
rect 9445 33768 9479 33802
rect 9445 33700 9479 33734
rect 7892 33576 7926 33610
rect 9445 33632 9479 33666
rect 7892 33508 7926 33542
rect 9445 33564 9479 33598
rect 9445 33496 9479 33530
rect 9667 34020 9701 34054
rect 9667 33952 9701 33986
rect 9667 33884 9701 33918
rect 9667 33816 9701 33850
rect 9667 33748 9701 33782
rect 9667 33680 9701 33714
rect 9667 33612 9701 33646
rect 9667 33544 9701 33578
rect 11525 34020 11559 34054
rect 11525 33952 11559 33986
rect 11525 33884 11559 33918
rect 11525 33816 11559 33850
rect 11525 33748 11559 33782
rect 11525 33680 11559 33714
rect 11525 33612 11559 33646
rect 11525 33544 11559 33578
rect 11747 34090 11781 34124
rect 11747 34022 11781 34056
rect 11747 33954 11781 33988
rect 11747 33886 11781 33920
rect 11747 33818 11781 33852
rect 11747 33750 11781 33784
rect 11747 33682 11781 33716
rect 11747 33614 11781 33648
rect 11747 33546 11781 33580
rect 7892 33440 7926 33474
rect 7892 33372 7926 33406
rect 7892 33304 7926 33338
rect 7052 33221 7086 33255
rect 7120 33221 7154 33255
rect 7188 33221 7222 33255
rect 7256 33221 7290 33255
rect 7324 33221 7358 33255
rect 7392 33221 7426 33255
rect 7460 33221 7494 33255
rect 7528 33221 7562 33255
rect 7596 33221 7630 33255
rect 7664 33221 7698 33255
rect 7732 33221 7766 33255
rect 7800 33221 7834 33255
rect 7868 33221 7902 33255
rect 9445 33428 9479 33462
rect 11747 33478 11781 33512
rect 11747 33410 11781 33444
rect 9445 33360 9479 33394
rect 9445 33292 9479 33326
rect 9445 33224 9479 33258
rect 11747 33342 11781 33376
rect 11747 33274 11781 33308
rect 9547 33200 9581 33234
rect 9615 33200 9649 33234
rect 9683 33200 9717 33234
rect 9751 33200 9785 33234
rect 9819 33200 9853 33234
rect 9887 33200 9921 33234
rect 9955 33200 9989 33234
rect 10023 33200 10057 33234
rect 10091 33200 10125 33234
rect 10159 33200 10193 33234
rect 10227 33200 10261 33234
rect 10295 33200 10329 33234
rect 10363 33200 10397 33234
rect 10431 33200 10465 33234
rect 10499 33200 10533 33234
rect 10567 33200 10601 33234
rect 10635 33200 10669 33234
rect 10703 33200 10737 33234
rect 10771 33200 10805 33234
rect 10839 33200 10873 33234
rect 10907 33200 10941 33234
rect 10975 33200 11009 33234
rect 11043 33200 11077 33234
rect 11111 33200 11145 33234
rect 11179 33200 11213 33234
rect 11247 33200 11281 33234
rect 11315 33200 11349 33234
rect 11383 33200 11417 33234
rect 11451 33200 11485 33234
rect 11519 33200 11553 33234
rect 11587 33200 11621 33234
rect 11655 33200 11689 33234
rect 11723 33200 11757 33234
rect 11877 34316 11911 34350
rect 11945 34316 11979 34350
rect 12013 34316 12047 34350
rect 12081 34316 12115 34350
rect 12149 34316 12183 34350
rect 12217 34316 12251 34350
rect 12285 34316 12319 34350
rect 12353 34316 12387 34350
rect 12421 34316 12455 34350
rect 12489 34316 12523 34350
rect 12557 34316 12591 34350
rect 12625 34316 12659 34350
rect 12693 34316 12727 34350
rect 12761 34316 12795 34350
rect 12885 34292 12919 34326
rect 11853 34207 11887 34241
rect 12002 34204 12036 34238
rect 12070 34204 12104 34238
rect 12138 34204 12172 34238
rect 12262 34204 12296 34238
rect 12330 34204 12364 34238
rect 12398 34204 12432 34238
rect 12505 34204 12539 34238
rect 12573 34204 12607 34238
rect 12641 34204 12675 34238
rect 12709 34204 12743 34238
rect 12885 34224 12919 34258
rect 11853 34139 11887 34173
rect 12885 34156 12919 34190
rect 11853 34071 11887 34105
rect 11853 34003 11887 34037
rect 11853 33935 11887 33969
rect 11853 33867 11887 33901
rect 11853 33799 11887 33833
rect 11853 33700 11887 33734
rect 11853 33632 11887 33666
rect 11853 33564 11887 33598
rect 11853 33496 11887 33530
rect 11853 33428 11887 33462
rect 12885 34088 12919 34122
rect 12885 34020 12919 34054
rect 12885 33952 12919 33986
rect 12885 33884 12919 33918
rect 12885 33816 12919 33850
rect 12885 33748 12919 33782
rect 12885 33680 12919 33714
rect 12885 33612 12919 33646
rect 12885 33544 12919 33578
rect 12885 33476 12919 33510
rect 11853 33360 11887 33394
rect 11853 33292 11887 33326
rect 12885 33408 12919 33442
rect 12885 33340 12919 33374
rect 11853 33224 11887 33258
rect 12885 33272 12919 33306
rect 11977 33200 12011 33234
rect 12045 33200 12079 33234
rect 12113 33200 12147 33234
rect 12181 33200 12215 33234
rect 12249 33200 12283 33234
rect 12317 33200 12351 33234
rect 12385 33200 12419 33234
rect 12453 33200 12487 33234
rect 12521 33200 12555 33234
rect 12589 33200 12623 33234
rect 12657 33200 12691 33234
rect 12725 33200 12759 33234
rect 12793 33200 12827 33234
rect 12861 33200 12895 33234
rect 13015 34317 13049 34351
rect 13083 34317 13117 34351
rect 13151 34317 13185 34351
rect 13219 34317 13253 34351
rect 13287 34317 13321 34351
rect 13355 34317 13389 34351
rect 13423 34317 13457 34351
rect 13491 34317 13525 34351
rect 13559 34317 13593 34351
rect 13627 34317 13661 34351
rect 13695 34317 13729 34351
rect 13763 34317 13797 34351
rect 13831 34317 13865 34351
rect 13899 34317 13933 34351
rect 13967 34317 14001 34351
rect 14035 34317 14069 34351
rect 14103 34317 14137 34351
rect 14171 34317 14205 34351
rect 14239 34317 14273 34351
rect 14307 34317 14341 34351
rect 14375 34317 14409 34351
rect 14443 34317 14477 34351
rect 14511 34317 14545 34351
rect 14579 34317 14613 34351
rect 14647 34317 14681 34351
rect 14715 34317 14749 34351
rect 14783 34317 14817 34351
rect 14851 34317 14885 34351
rect 14919 34317 14953 34351
rect 14987 34317 15021 34351
rect 15055 34317 15089 34351
rect 15123 34317 15157 34351
rect 15227 34318 15261 34352
rect 15295 34318 15329 34352
rect 15363 34318 15397 34352
rect 15431 34318 15465 34352
rect 15499 34318 15533 34352
rect 15567 34318 15601 34352
rect 15635 34318 15669 34352
rect 15703 34318 15737 34352
rect 15771 34318 15805 34352
rect 15839 34318 15873 34352
rect 15907 34318 15941 34352
rect 15975 34318 16009 34352
rect 16043 34318 16077 34352
rect 12991 34244 13025 34278
rect 16159 34294 16193 34328
rect 12991 34176 13025 34210
rect 13119 34186 13153 34220
rect 13187 34186 13221 34220
rect 13255 34186 13289 34220
rect 13323 34186 13357 34220
rect 13391 34186 13425 34220
rect 13459 34186 13493 34220
rect 13527 34186 13561 34220
rect 13595 34186 13629 34220
rect 13663 34186 13697 34220
rect 13731 34186 13765 34220
rect 13893 34186 13927 34220
rect 13961 34186 13995 34220
rect 14029 34186 14063 34220
rect 14097 34186 14131 34220
rect 14165 34186 14199 34220
rect 14233 34186 14267 34220
rect 14301 34186 14335 34220
rect 14369 34186 14403 34220
rect 14437 34186 14471 34220
rect 14505 34186 14539 34220
rect 16159 34226 16193 34260
rect 12991 34108 13025 34142
rect 16159 34158 16193 34192
rect 12991 34040 13025 34074
rect 12991 33972 13025 34006
rect 12991 33904 13025 33938
rect 12991 33836 13025 33870
rect 12991 33768 13025 33802
rect 12991 33700 13025 33734
rect 12991 33632 13025 33666
rect 12991 33564 13025 33598
rect 12991 33496 13025 33530
rect 12991 33428 13025 33462
rect 16159 34090 16193 34124
rect 16159 34022 16193 34056
rect 16159 33954 16193 33988
rect 16159 33886 16193 33920
rect 16159 33818 16193 33852
rect 16159 33750 16193 33784
rect 16159 33682 16193 33716
rect 16159 33614 16193 33648
rect 16159 33546 16193 33580
rect 16159 33478 16193 33512
rect 12991 33360 13025 33394
rect 16159 33410 16193 33444
rect 16159 33342 16193 33376
rect 12991 33292 13025 33326
rect 12991 33224 13025 33258
rect 16159 33274 16193 33308
rect 13106 33200 13140 33234
rect 13174 33200 13208 33234
rect 13242 33200 13276 33234
rect 13310 33200 13344 33234
rect 13378 33200 13412 33234
rect 13446 33200 13480 33234
rect 13514 33200 13548 33234
rect 13582 33200 13616 33234
rect 13650 33200 13684 33234
rect 13718 33200 13752 33234
rect 13786 33200 13820 33234
rect 13854 33200 13888 33234
rect 13922 33200 13956 33234
rect 13990 33200 14024 33234
rect 14058 33200 14092 33234
rect 14126 33200 14160 33234
rect 14194 33200 14228 33234
rect 14262 33200 14296 33234
rect 14330 33200 14364 33234
rect 14398 33200 14432 33234
rect 14466 33200 14500 33234
rect 14534 33200 14568 33234
rect 14639 33200 14673 33234
rect 14707 33200 14741 33234
rect 14775 33200 14809 33234
rect 14843 33200 14877 33234
rect 14911 33200 14945 33234
rect 14979 33200 15013 33234
rect 15047 33200 15081 33234
rect 15115 33200 15149 33234
rect 15183 33200 15217 33234
rect 15251 33200 15285 33234
rect 15319 33200 15353 33234
rect 15387 33200 15421 33234
rect 15455 33200 15489 33234
rect 15523 33200 15557 33234
rect 15591 33200 15625 33234
rect 15659 33200 15693 33234
rect 15727 33200 15761 33234
rect 15795 33200 15829 33234
rect 15863 33200 15897 33234
rect 15931 33200 15965 33234
rect 15999 33200 16033 33234
rect 16067 33200 16101 33234
rect 16135 33200 16169 33234
rect 11481 19226 11515 19260
rect 11549 19226 11583 19260
rect 11617 19226 11651 19260
rect 11685 19226 11719 19260
rect 11753 19226 11787 19260
rect 11821 19226 11855 19260
rect 11889 19226 11923 19260
rect 11957 19226 11991 19260
rect 12025 19226 12059 19260
rect 12093 19226 12127 19260
rect 12161 19226 12195 19260
rect 12229 19226 12263 19260
rect 12297 19226 12331 19260
rect 12365 19226 12399 19260
rect 12433 19226 12467 19260
rect 12501 19226 12535 19260
rect 12569 19226 12603 19260
rect 12637 19226 12671 19260
rect 12705 19226 12739 19260
rect 12773 19226 12807 19260
rect 12841 19226 12875 19260
rect 12909 19226 12943 19260
rect 12977 19226 13011 19260
rect 13045 19226 13079 19260
rect 13113 19226 13147 19260
rect 13181 19226 13215 19260
rect 13249 19226 13283 19260
rect 13317 19226 13351 19260
rect 13385 19226 13419 19260
rect 13453 19226 13487 19260
rect 13521 19226 13555 19260
rect 13589 19226 13623 19260
rect 13657 19226 13691 19260
rect 13725 19226 13759 19260
rect 13793 19226 13827 19260
rect 13861 19226 13895 19260
rect 13929 19226 13963 19260
rect 13997 19226 14031 19260
rect 14065 19226 14099 19260
rect 14133 19226 14167 19260
rect 14201 19226 14235 19260
rect 14269 19226 14303 19260
rect 14360 19226 14394 19260
rect 14428 19226 14462 19260
rect 14496 19226 14530 19260
rect 14564 19226 14598 19260
rect 14632 19226 14666 19260
rect 14700 19226 14734 19260
rect 14768 19226 14802 19260
rect 14836 19226 14870 19260
rect 14904 19226 14938 19260
rect 14972 19226 15006 19260
rect 15040 19226 15074 19260
rect 15108 19226 15142 19260
rect 15176 19226 15210 19260
rect 15244 19226 15278 19260
rect 15312 19226 15346 19260
rect 15380 19226 15414 19260
rect 15448 19226 15482 19260
rect 15516 19226 15550 19260
rect 15584 19226 15618 19260
rect 15652 19226 15686 19260
rect 15720 19226 15754 19260
rect 15788 19226 15822 19260
rect 15856 19226 15890 19260
rect 15924 19226 15958 19260
rect 15992 19226 16026 19260
rect 16060 19226 16094 19260
rect 16128 19226 16162 19260
rect 16196 19226 16230 19260
rect 16264 19226 16298 19260
rect 16332 19226 16366 19260
rect 16400 19226 16434 19260
rect 16468 19226 16502 19260
rect 16536 19226 16570 19260
rect 16604 19226 16638 19260
rect 16672 19226 16706 19260
rect 16740 19226 16774 19260
rect 16808 19226 16842 19260
rect 16876 19226 16910 19260
rect 16944 19226 16978 19260
rect 17012 19226 17046 19260
rect 17080 19226 17114 19260
rect 11457 19132 11491 19166
rect 11457 19064 11491 19098
rect 11457 18996 11491 19030
rect 11457 18928 11491 18962
rect 11457 18860 11491 18894
rect 11457 18792 11491 18826
rect 11457 18724 11491 18758
rect 11457 18656 11491 18690
rect 11457 18588 11491 18622
rect 11457 18520 11491 18554
rect 11457 18452 11491 18486
rect 11457 18384 11491 18418
rect 11457 18316 11491 18350
rect 11457 18248 11491 18282
rect 11457 18180 11491 18214
rect 11457 18112 11491 18146
rect 11457 18044 11491 18078
rect 11457 17976 11491 18010
rect 11457 17908 11491 17942
rect 11457 17840 11491 17874
rect 11457 17772 11491 17806
rect 11457 17704 11491 17738
rect 11457 17636 11491 17670
rect 17181 19202 17215 19236
rect 17181 19134 17215 19168
rect 17181 19066 17215 19100
rect 17181 18998 17215 19032
rect 17181 18930 17215 18964
rect 17181 18862 17215 18896
rect 17181 18794 17215 18828
rect 17181 18726 17215 18760
rect 17181 18658 17215 18692
rect 17181 18590 17215 18624
rect 17181 18522 17215 18556
rect 17181 18454 17215 18488
rect 17181 18386 17215 18420
rect 17181 18318 17215 18352
rect 17181 18250 17215 18284
rect 17181 18182 17215 18216
rect 17181 18114 17215 18148
rect 17181 18046 17215 18080
rect 17181 17978 17215 18012
rect 17181 17910 17215 17944
rect 17181 17842 17215 17876
rect 17181 17774 17215 17808
rect 17181 17706 17215 17740
rect 17181 17638 17215 17672
rect 11457 17568 11491 17602
rect 11457 17500 11491 17534
rect 11457 17432 11491 17466
rect 11457 17364 11491 17398
rect 11457 17296 11491 17330
rect 11457 17228 11491 17262
rect 11457 17160 11491 17194
rect 11457 17092 11491 17126
rect 11457 17024 11491 17058
rect 11457 16956 11491 16990
rect 11457 16888 11491 16922
rect 11457 16820 11491 16854
rect 11457 16752 11491 16786
rect 11457 16684 11491 16718
rect 11457 16616 11491 16650
rect 11457 16548 11491 16582
rect 11457 16480 11491 16514
rect 11457 16412 11491 16446
rect 8988 16312 9022 16346
rect 9056 16312 9090 16346
rect 9124 16312 9158 16346
rect 9192 16312 9226 16346
rect 9260 16312 9294 16346
rect 9328 16312 9362 16346
rect 9396 16312 9430 16346
rect 9464 16312 9498 16346
rect 9532 16312 9566 16346
rect 9600 16312 9634 16346
rect 9668 16312 9702 16346
rect 9736 16312 9770 16346
rect 9804 16312 9838 16346
rect 8964 16232 8998 16266
rect 8964 16164 8998 16198
rect 8964 16096 8998 16130
rect 8964 16028 8998 16062
rect 8964 15960 8998 15994
rect 8964 15892 8998 15926
rect 8964 15824 8998 15858
rect 8964 15756 8998 15790
rect 8964 15688 8998 15722
rect 8964 15620 8998 15654
rect 8964 15481 8998 15515
rect 8964 15413 8998 15447
rect 8964 15345 8998 15379
rect 8964 15277 8998 15311
rect 8964 15209 8998 15243
rect 8964 15141 8998 15175
rect 8964 15073 8998 15107
rect 8964 15005 8998 15039
rect 8964 14937 8998 14971
rect 8964 14869 8998 14903
rect 9904 16288 9938 16322
rect 9904 16220 9938 16254
rect 9904 16152 9938 16186
rect 9904 16084 9938 16118
rect 9904 16016 9938 16050
rect 11457 16344 11491 16378
rect 11457 16276 11491 16310
rect 11457 16208 11491 16242
rect 11457 16140 11491 16174
rect 11457 16072 11491 16106
rect 17181 17570 17215 17604
rect 17181 17502 17215 17536
rect 17181 17434 17215 17468
rect 17181 17366 17215 17400
rect 17181 17298 17215 17332
rect 17181 17230 17215 17264
rect 17181 17162 17215 17196
rect 17181 17094 17215 17128
rect 17181 17026 17215 17060
rect 17181 16958 17215 16992
rect 17181 16890 17215 16924
rect 17181 16822 17215 16856
rect 17181 16754 17215 16788
rect 17181 16686 17215 16720
rect 17181 16618 17215 16652
rect 17181 16550 17215 16584
rect 17181 16482 17215 16516
rect 17181 16414 17215 16448
rect 17181 16346 17215 16380
rect 17181 16278 17215 16312
rect 17181 16210 17215 16244
rect 17181 16142 17215 16176
rect 11581 16048 11615 16082
rect 11649 16048 11683 16082
rect 11717 16048 11751 16082
rect 11785 16048 11819 16082
rect 11853 16048 11887 16082
rect 11921 16048 11955 16082
rect 11989 16048 12023 16082
rect 12057 16048 12091 16082
rect 12125 16048 12159 16082
rect 12193 16048 12227 16082
rect 12261 16048 12295 16082
rect 12329 16048 12363 16082
rect 12397 16048 12431 16082
rect 12465 16048 12499 16082
rect 12533 16048 12567 16082
rect 12601 16048 12635 16082
rect 12669 16048 12703 16082
rect 12737 16048 12771 16082
rect 12805 16048 12839 16082
rect 12873 16048 12907 16082
rect 12941 16048 12975 16082
rect 13009 16048 13043 16082
rect 13077 16048 13111 16082
rect 13145 16048 13179 16082
rect 13213 16048 13247 16082
rect 13281 16048 13315 16082
rect 13349 16048 13383 16082
rect 13417 16048 13451 16082
rect 13485 16048 13519 16082
rect 13553 16048 13587 16082
rect 13621 16048 13655 16082
rect 13689 16048 13723 16082
rect 13757 16048 13791 16082
rect 13825 16048 13859 16082
rect 13893 16048 13927 16082
rect 13961 16048 13995 16082
rect 14029 16048 14063 16082
rect 14097 16048 14131 16082
rect 14165 16048 14199 16082
rect 14233 16048 14267 16082
rect 14301 16048 14335 16082
rect 14369 16048 14403 16082
rect 14437 16048 14471 16082
rect 14505 16048 14539 16082
rect 14573 16048 14607 16082
rect 14641 16048 14675 16082
rect 14709 16048 14743 16082
rect 14777 16048 14811 16082
rect 14845 16048 14879 16082
rect 14913 16048 14947 16082
rect 14981 16048 15015 16082
rect 15049 16048 15083 16082
rect 15117 16048 15151 16082
rect 15185 16048 15219 16082
rect 15253 16048 15287 16082
rect 15321 16048 15355 16082
rect 15389 16048 15423 16082
rect 15457 16048 15491 16082
rect 15525 16048 15559 16082
rect 15593 16048 15627 16082
rect 15661 16048 15695 16082
rect 15729 16048 15763 16082
rect 15797 16048 15831 16082
rect 15865 16048 15899 16082
rect 15933 16048 15967 16082
rect 16001 16048 16035 16082
rect 16069 16048 16103 16082
rect 16137 16048 16171 16082
rect 16205 16048 16239 16082
rect 16273 16048 16307 16082
rect 16341 16048 16375 16082
rect 16409 16048 16443 16082
rect 16477 16048 16511 16082
rect 16545 16048 16579 16082
rect 16613 16048 16647 16082
rect 16681 16048 16715 16082
rect 16749 16048 16783 16082
rect 16817 16048 16851 16082
rect 16885 16048 16919 16082
rect 16953 16048 16987 16082
rect 17021 16048 17055 16082
rect 17089 16048 17123 16082
rect 17157 16048 17191 16082
rect 17287 19202 17321 19236
rect 17383 19226 17417 19260
rect 17451 19226 17485 19260
rect 17519 19226 17553 19260
rect 17587 19226 17621 19260
rect 17655 19226 17689 19260
rect 17723 19226 17757 19260
rect 17791 19226 17825 19260
rect 17859 19226 17893 19260
rect 17927 19226 17961 19260
rect 17995 19226 18029 19260
rect 18063 19226 18097 19260
rect 18131 19226 18165 19260
rect 18199 19226 18233 19260
rect 18267 19226 18301 19260
rect 18335 19226 18369 19260
rect 18403 19226 18437 19260
rect 18471 19226 18505 19260
rect 18539 19226 18573 19260
rect 18607 19226 18641 19260
rect 18675 19226 18709 19260
rect 18743 19226 18777 19260
rect 18811 19226 18845 19260
rect 18879 19226 18913 19260
rect 18947 19226 18981 19260
rect 19015 19226 19049 19260
rect 19083 19226 19117 19260
rect 19151 19226 19185 19260
rect 19219 19226 19253 19260
rect 19287 19226 19321 19260
rect 19355 19226 19389 19260
rect 19423 19226 19457 19260
rect 19491 19226 19525 19260
rect 19559 19226 19593 19260
rect 19627 19226 19661 19260
rect 19695 19226 19729 19260
rect 19763 19226 19797 19260
rect 19831 19226 19865 19260
rect 19899 19226 19933 19260
rect 19967 19226 20001 19260
rect 20035 19226 20069 19260
rect 20103 19226 20137 19260
rect 20171 19226 20205 19260
rect 17287 19134 17321 19168
rect 17287 19066 17321 19100
rect 17287 18998 17321 19032
rect 17287 18930 17321 18964
rect 17287 18862 17321 18896
rect 17287 18794 17321 18828
rect 17287 18726 17321 18760
rect 17287 18658 17321 18692
rect 17287 18590 17321 18624
rect 17287 18522 17321 18556
rect 17287 18454 17321 18488
rect 17287 18386 17321 18420
rect 17287 18318 17321 18352
rect 17287 18250 17321 18284
rect 17287 18182 17321 18216
rect 17287 18114 17321 18148
rect 17287 18046 17321 18080
rect 17287 17978 17321 18012
rect 17287 17910 17321 17944
rect 17287 17842 17321 17876
rect 17287 17774 17321 17808
rect 17287 17706 17321 17740
rect 17287 17638 17321 17672
rect 17287 17570 17321 17604
rect 17287 17502 17321 17536
rect 17287 17434 17321 17468
rect 17287 17366 17321 17400
rect 17287 17298 17321 17332
rect 17287 17230 17321 17264
rect 17287 17162 17321 17196
rect 17287 17094 17321 17128
rect 17287 17026 17321 17060
rect 17287 16958 17321 16992
rect 17287 16890 17321 16924
rect 17287 16822 17321 16856
rect 17287 16754 17321 16788
rect 17287 16686 17321 16720
rect 17287 16618 17321 16652
rect 17287 16550 17321 16584
rect 17287 16482 17321 16516
rect 17287 16414 17321 16448
rect 17287 16346 17321 16380
rect 17287 16278 17321 16312
rect 17287 16210 17321 16244
rect 17287 16142 17321 16176
rect 20195 19106 20229 19140
rect 20195 19038 20229 19072
rect 20195 18970 20229 19004
rect 20195 18902 20229 18936
rect 20195 18834 20229 18868
rect 20195 18766 20229 18800
rect 20195 18698 20229 18732
rect 20195 18630 20229 18664
rect 20195 18562 20229 18596
rect 20195 18494 20229 18528
rect 20195 18426 20229 18460
rect 20195 18358 20229 18392
rect 20195 18290 20229 18324
rect 20195 18222 20229 18256
rect 20195 18154 20229 18188
rect 20195 18086 20229 18120
rect 20195 18018 20229 18052
rect 20195 17950 20229 17984
rect 20195 17882 20229 17916
rect 20195 17814 20229 17848
rect 20195 17746 20229 17780
rect 20195 17678 20229 17712
rect 20195 17568 20229 17602
rect 20195 17500 20229 17534
rect 20195 17432 20229 17466
rect 20195 17364 20229 17398
rect 20195 17296 20229 17330
rect 20195 17228 20229 17262
rect 20195 17160 20229 17194
rect 20195 17092 20229 17126
rect 20195 17024 20229 17058
rect 20195 16956 20229 16990
rect 20195 16888 20229 16922
rect 20195 16820 20229 16854
rect 20195 16752 20229 16786
rect 20195 16684 20229 16718
rect 20195 16616 20229 16650
rect 20195 16548 20229 16582
rect 20195 16480 20229 16514
rect 20195 16412 20229 16446
rect 20195 16344 20229 16378
rect 20195 16276 20229 16310
rect 20195 16208 20229 16242
rect 20195 16140 20229 16174
rect 17311 16048 17345 16082
rect 17379 16048 17413 16082
rect 17447 16048 17481 16082
rect 17515 16048 17549 16082
rect 17583 16048 17617 16082
rect 17651 16048 17685 16082
rect 17719 16048 17753 16082
rect 17787 16048 17821 16082
rect 17855 16048 17889 16082
rect 17923 16048 17957 16082
rect 17991 16048 18025 16082
rect 18059 16048 18093 16082
rect 18127 16048 18161 16082
rect 18195 16048 18229 16082
rect 18263 16048 18297 16082
rect 18331 16048 18365 16082
rect 18399 16048 18433 16082
rect 18467 16048 18501 16082
rect 18535 16048 18569 16082
rect 18603 16048 18637 16082
rect 18671 16048 18705 16082
rect 18739 16048 18773 16082
rect 18807 16048 18841 16082
rect 18875 16048 18909 16082
rect 18943 16048 18977 16082
rect 19011 16048 19045 16082
rect 19079 16048 19113 16082
rect 19147 16048 19181 16082
rect 19215 16048 19249 16082
rect 19283 16048 19317 16082
rect 19351 16048 19385 16082
rect 19419 16048 19453 16082
rect 19487 16048 19521 16082
rect 19555 16048 19589 16082
rect 19623 16048 19657 16082
rect 19691 16048 19725 16082
rect 19759 16048 19793 16082
rect 19827 16048 19861 16082
rect 19895 16048 19929 16082
rect 19963 16048 19997 16082
rect 20031 16048 20065 16082
rect 20099 16048 20133 16082
rect 20195 16072 20229 16106
rect 20301 19202 20335 19236
rect 20374 19226 20408 19260
rect 20442 19226 20476 19260
rect 20510 19226 20544 19260
rect 20578 19226 20612 19260
rect 20646 19226 20680 19260
rect 20714 19226 20748 19260
rect 20782 19226 20816 19260
rect 20850 19226 20884 19260
rect 20918 19226 20952 19260
rect 20986 19226 21020 19260
rect 21054 19226 21088 19260
rect 21122 19226 21156 19260
rect 21190 19226 21224 19260
rect 21258 19226 21292 19260
rect 21326 19226 21360 19260
rect 21394 19226 21428 19260
rect 21462 19226 21496 19260
rect 21530 19226 21564 19260
rect 21598 19226 21632 19260
rect 21666 19226 21700 19260
rect 21734 19226 21768 19260
rect 21802 19226 21836 19260
rect 21870 19226 21904 19260
rect 21938 19226 21972 19260
rect 22006 19226 22040 19260
rect 22074 19226 22108 19260
rect 22142 19226 22176 19260
rect 22210 19226 22244 19260
rect 22278 19226 22312 19260
rect 22346 19226 22380 19260
rect 22414 19226 22448 19260
rect 22482 19226 22516 19260
rect 22550 19226 22584 19260
rect 22618 19226 22652 19260
rect 22686 19226 22720 19260
rect 22754 19226 22788 19260
rect 22822 19226 22856 19260
rect 22890 19226 22924 19260
rect 22958 19226 22992 19260
rect 23026 19226 23060 19260
rect 23157 19226 23191 19260
rect 23225 19226 23259 19260
rect 23293 19226 23327 19260
rect 23361 19226 23395 19260
rect 23429 19226 23463 19260
rect 23497 19226 23531 19260
rect 23565 19226 23599 19260
rect 23633 19226 23667 19260
rect 23701 19226 23735 19260
rect 23769 19226 23803 19260
rect 23837 19226 23871 19260
rect 23905 19226 23939 19260
rect 23973 19226 24007 19260
rect 24041 19226 24075 19260
rect 24109 19226 24143 19260
rect 24177 19226 24211 19260
rect 24245 19226 24279 19260
rect 24313 19226 24347 19260
rect 24381 19226 24415 19260
rect 24449 19226 24483 19260
rect 24517 19226 24551 19260
rect 24585 19226 24619 19260
rect 24653 19226 24687 19260
rect 24721 19226 24755 19260
rect 24789 19226 24823 19260
rect 24857 19226 24891 19260
rect 24925 19226 24959 19260
rect 24993 19226 25027 19260
rect 25061 19226 25095 19260
rect 25129 19226 25163 19260
rect 25197 19226 25231 19260
rect 25265 19226 25299 19260
rect 25333 19226 25367 19260
rect 25401 19226 25435 19260
rect 25469 19226 25503 19260
rect 25537 19226 25571 19260
rect 25605 19226 25639 19260
rect 25673 19226 25707 19260
rect 25741 19226 25775 19260
rect 25809 19226 25843 19260
rect 20301 19134 20335 19168
rect 20301 19066 20335 19100
rect 20301 18998 20335 19032
rect 20301 18930 20335 18964
rect 20301 18862 20335 18896
rect 20301 18794 20335 18828
rect 20301 18726 20335 18760
rect 20301 18658 20335 18692
rect 20301 18590 20335 18624
rect 20301 18522 20335 18556
rect 20301 18454 20335 18488
rect 20301 18386 20335 18420
rect 20301 18318 20335 18352
rect 20301 18250 20335 18284
rect 20301 18182 20335 18216
rect 20301 18114 20335 18148
rect 20301 18046 20335 18080
rect 20301 17978 20335 18012
rect 20301 17910 20335 17944
rect 20301 17842 20335 17876
rect 20301 17774 20335 17808
rect 20301 17706 20335 17740
rect 20301 17638 20335 17672
rect 20301 17570 20335 17604
rect 20301 17502 20335 17536
rect 20301 17434 20335 17468
rect 20301 17366 20335 17400
rect 20301 17298 20335 17332
rect 20301 17230 20335 17264
rect 20301 17162 20335 17196
rect 20301 17094 20335 17128
rect 20301 17026 20335 17060
rect 20301 16958 20335 16992
rect 20301 16890 20335 16924
rect 20301 16822 20335 16856
rect 20301 16754 20335 16788
rect 20301 16686 20335 16720
rect 20301 16618 20335 16652
rect 20301 16550 20335 16584
rect 20301 16482 20335 16516
rect 20301 16414 20335 16448
rect 20301 16346 20335 16380
rect 20301 16278 20335 16312
rect 20301 16210 20335 16244
rect 20301 16142 20335 16176
rect 25833 19132 25867 19166
rect 25833 19064 25867 19098
rect 25833 18996 25867 19030
rect 25833 18928 25867 18962
rect 25833 18860 25867 18894
rect 25833 18792 25867 18826
rect 25833 18724 25867 18758
rect 25833 18656 25867 18690
rect 25833 18588 25867 18622
rect 25833 18520 25867 18554
rect 25833 18452 25867 18486
rect 25833 18384 25867 18418
rect 25833 18316 25867 18350
rect 25833 18248 25867 18282
rect 25833 18180 25867 18214
rect 25833 18112 25867 18146
rect 25833 18044 25867 18078
rect 25833 17976 25867 18010
rect 25833 17908 25867 17942
rect 25833 17840 25867 17874
rect 25833 17772 25867 17806
rect 25833 17704 25867 17738
rect 25833 17636 25867 17670
rect 25833 17568 25867 17602
rect 25833 17500 25867 17534
rect 25833 17432 25867 17466
rect 25833 17364 25867 17398
rect 25833 17296 25867 17330
rect 25833 17228 25867 17262
rect 25833 17160 25867 17194
rect 25833 17092 25867 17126
rect 25833 17024 25867 17058
rect 25833 16956 25867 16990
rect 25833 16888 25867 16922
rect 25833 16820 25867 16854
rect 25833 16752 25867 16786
rect 25833 16684 25867 16718
rect 25833 16616 25867 16650
rect 25833 16548 25867 16582
rect 25833 16480 25867 16514
rect 25833 16412 25867 16446
rect 25833 16344 25867 16378
rect 25833 16276 25867 16310
rect 25833 16208 25867 16242
rect 25833 16140 25867 16174
rect 20325 16048 20359 16082
rect 20393 16048 20427 16082
rect 20461 16048 20495 16082
rect 20529 16048 20563 16082
rect 20597 16048 20631 16082
rect 20665 16048 20699 16082
rect 20733 16048 20767 16082
rect 20801 16048 20835 16082
rect 20869 16048 20903 16082
rect 20937 16048 20971 16082
rect 21005 16048 21039 16082
rect 21073 16048 21107 16082
rect 21141 16048 21175 16082
rect 21209 16048 21243 16082
rect 21277 16048 21311 16082
rect 21345 16048 21379 16082
rect 21413 16048 21447 16082
rect 21481 16048 21515 16082
rect 21549 16048 21583 16082
rect 21617 16048 21651 16082
rect 21685 16048 21719 16082
rect 21753 16048 21787 16082
rect 21821 16048 21855 16082
rect 21889 16048 21923 16082
rect 21957 16048 21991 16082
rect 22025 16048 22059 16082
rect 22093 16048 22127 16082
rect 22161 16048 22195 16082
rect 22229 16048 22263 16082
rect 22297 16048 22331 16082
rect 22365 16048 22399 16082
rect 22433 16048 22467 16082
rect 22501 16048 22535 16082
rect 22569 16048 22603 16082
rect 22637 16048 22671 16082
rect 22705 16048 22739 16082
rect 22773 16048 22807 16082
rect 22841 16048 22875 16082
rect 22909 16048 22943 16082
rect 22977 16048 23011 16082
rect 23045 16048 23079 16082
rect 23113 16048 23147 16082
rect 23181 16048 23215 16082
rect 23249 16048 23283 16082
rect 23317 16048 23351 16082
rect 23385 16048 23419 16082
rect 23453 16048 23487 16082
rect 23521 16048 23555 16082
rect 23589 16048 23623 16082
rect 23657 16048 23691 16082
rect 23725 16048 23759 16082
rect 23793 16048 23827 16082
rect 23861 16048 23895 16082
rect 23929 16048 23963 16082
rect 23997 16048 24031 16082
rect 24065 16048 24099 16082
rect 24133 16048 24167 16082
rect 24201 16048 24235 16082
rect 24269 16048 24303 16082
rect 24337 16048 24371 16082
rect 24405 16048 24439 16082
rect 24473 16048 24507 16082
rect 24541 16048 24575 16082
rect 24609 16048 24643 16082
rect 24677 16048 24711 16082
rect 24745 16048 24779 16082
rect 24813 16048 24847 16082
rect 24881 16048 24915 16082
rect 24949 16048 24983 16082
rect 25017 16048 25051 16082
rect 25085 16048 25119 16082
rect 25153 16048 25187 16082
rect 25221 16048 25255 16082
rect 25289 16048 25323 16082
rect 25357 16048 25391 16082
rect 25425 16048 25459 16082
rect 25493 16048 25527 16082
rect 25561 16048 25595 16082
rect 25629 16048 25663 16082
rect 25697 16048 25731 16082
rect 25765 16048 25799 16082
rect 25833 16072 25867 16106
rect 9904 15948 9938 15982
rect 9904 15880 9938 15914
rect 9904 15812 9938 15846
rect 9904 15744 9938 15778
rect 9904 15676 9938 15710
rect 9904 15608 9938 15642
rect 9904 15540 9938 15574
rect 9904 15472 9938 15506
rect 9904 15404 9938 15438
rect 9904 15336 9938 15370
rect 9904 15268 9938 15302
rect 11481 15942 11515 15976
rect 11549 15942 11583 15976
rect 11617 15942 11651 15976
rect 11685 15942 11719 15976
rect 11753 15942 11787 15976
rect 11821 15942 11855 15976
rect 11889 15942 11923 15976
rect 11957 15942 11991 15976
rect 12025 15942 12059 15976
rect 12093 15942 12127 15976
rect 12161 15942 12195 15976
rect 12229 15942 12263 15976
rect 12297 15942 12331 15976
rect 12365 15942 12399 15976
rect 12433 15942 12467 15976
rect 12501 15942 12535 15976
rect 12649 15942 12683 15976
rect 12717 15942 12751 15976
rect 12785 15942 12819 15976
rect 12853 15942 12887 15976
rect 12921 15942 12955 15976
rect 12989 15942 13023 15976
rect 13057 15942 13091 15976
rect 13125 15942 13159 15976
rect 13193 15942 13227 15976
rect 13261 15942 13295 15976
rect 13329 15942 13363 15976
rect 13397 15942 13431 15976
rect 13465 15942 13499 15976
rect 13533 15942 13567 15976
rect 13601 15942 13635 15976
rect 13669 15942 13703 15976
rect 11457 15868 11491 15902
rect 11457 15800 11491 15834
rect 11457 15732 11491 15766
rect 11457 15664 11491 15698
rect 11457 15596 11491 15630
rect 11457 15528 11491 15562
rect 11457 15460 11491 15494
rect 11457 15392 11491 15426
rect 11457 15324 11491 15358
rect 9904 15200 9938 15234
rect 11457 15256 11491 15290
rect 9904 15132 9938 15166
rect 11457 15188 11491 15222
rect 11457 15120 11491 15154
rect 9904 15064 9938 15098
rect 9904 14996 9938 15030
rect 9904 14928 9938 14962
rect 9064 14845 9098 14879
rect 9132 14845 9166 14879
rect 9200 14845 9234 14879
rect 9268 14845 9302 14879
rect 9336 14845 9370 14879
rect 9404 14845 9438 14879
rect 9472 14845 9506 14879
rect 9540 14845 9574 14879
rect 9608 14845 9642 14879
rect 9676 14845 9710 14879
rect 9744 14845 9778 14879
rect 9812 14845 9846 14879
rect 9880 14845 9914 14879
rect 11457 15052 11491 15086
rect 11457 14984 11491 15018
rect 11457 14916 11491 14950
rect 11457 14848 11491 14882
rect 13759 15918 13793 15952
rect 13759 15850 13793 15884
rect 13759 15782 13793 15816
rect 13759 15714 13793 15748
rect 13759 15646 13793 15680
rect 13759 15578 13793 15612
rect 13759 15510 13793 15544
rect 13759 15442 13793 15476
rect 13759 15374 13793 15408
rect 13759 15306 13793 15340
rect 13759 15238 13793 15272
rect 13759 15170 13793 15204
rect 13759 15102 13793 15136
rect 13759 15034 13793 15068
rect 13759 14966 13793 15000
rect 13759 14898 13793 14932
rect 11559 14824 11593 14858
rect 11627 14824 11661 14858
rect 11695 14824 11729 14858
rect 11763 14824 11797 14858
rect 11831 14824 11865 14858
rect 11899 14824 11933 14858
rect 11967 14824 12001 14858
rect 12035 14824 12069 14858
rect 12103 14824 12137 14858
rect 12171 14824 12205 14858
rect 12239 14824 12273 14858
rect 12307 14824 12341 14858
rect 12375 14824 12409 14858
rect 12443 14824 12477 14858
rect 12511 14824 12545 14858
rect 12579 14824 12613 14858
rect 12647 14824 12681 14858
rect 12715 14824 12749 14858
rect 12783 14824 12817 14858
rect 12851 14824 12885 14858
rect 12919 14824 12953 14858
rect 12987 14824 13021 14858
rect 13055 14824 13089 14858
rect 13123 14824 13157 14858
rect 13191 14824 13225 14858
rect 13259 14824 13293 14858
rect 13327 14824 13361 14858
rect 13395 14824 13429 14858
rect 13463 14824 13497 14858
rect 13531 14824 13565 14858
rect 13599 14824 13633 14858
rect 13667 14824 13701 14858
rect 13735 14824 13769 14858
rect 13889 15940 13923 15974
rect 13957 15940 13991 15974
rect 14025 15940 14059 15974
rect 14093 15940 14127 15974
rect 14161 15940 14195 15974
rect 14229 15940 14263 15974
rect 14297 15940 14331 15974
rect 14365 15940 14399 15974
rect 14433 15940 14467 15974
rect 14501 15940 14535 15974
rect 14569 15940 14603 15974
rect 14637 15940 14671 15974
rect 14705 15940 14739 15974
rect 14773 15940 14807 15974
rect 13865 15831 13899 15865
rect 13865 15763 13899 15797
rect 13865 15695 13899 15729
rect 13865 15627 13899 15661
rect 13865 15559 13899 15593
rect 13865 15491 13899 15525
rect 13865 15423 13899 15457
rect 13865 15324 13899 15358
rect 13865 15256 13899 15290
rect 13865 15188 13899 15222
rect 13865 15120 13899 15154
rect 13865 15052 13899 15086
rect 13865 14984 13899 15018
rect 13865 14916 13899 14950
rect 13865 14848 13899 14882
rect 14897 15916 14931 15950
rect 14897 15848 14931 15882
rect 14897 15780 14931 15814
rect 14897 15712 14931 15746
rect 14897 15644 14931 15678
rect 14897 15576 14931 15610
rect 14897 15508 14931 15542
rect 14897 15440 14931 15474
rect 14897 15372 14931 15406
rect 14897 15304 14931 15338
rect 14897 15236 14931 15270
rect 14897 15168 14931 15202
rect 14897 15100 14931 15134
rect 14897 15032 14931 15066
rect 14897 14964 14931 14998
rect 14897 14896 14931 14930
rect 13989 14824 14023 14858
rect 14057 14824 14091 14858
rect 14125 14824 14159 14858
rect 14193 14824 14227 14858
rect 14261 14824 14295 14858
rect 14329 14824 14363 14858
rect 14397 14824 14431 14858
rect 14465 14824 14499 14858
rect 14533 14824 14567 14858
rect 14601 14824 14635 14858
rect 14669 14824 14703 14858
rect 14737 14824 14771 14858
rect 14805 14824 14839 14858
rect 14873 14824 14907 14858
rect 15027 15941 15061 15975
rect 15095 15941 15129 15975
rect 15163 15941 15197 15975
rect 15231 15941 15265 15975
rect 15299 15941 15333 15975
rect 15367 15941 15401 15975
rect 15435 15941 15469 15975
rect 15503 15941 15537 15975
rect 15571 15941 15605 15975
rect 15639 15941 15673 15975
rect 15707 15941 15741 15975
rect 15775 15941 15809 15975
rect 15843 15941 15877 15975
rect 15911 15941 15945 15975
rect 15979 15941 16013 15975
rect 16047 15941 16081 15975
rect 16115 15941 16149 15975
rect 16183 15941 16217 15975
rect 16251 15941 16285 15975
rect 16319 15941 16353 15975
rect 16387 15941 16421 15975
rect 16455 15941 16489 15975
rect 16523 15941 16557 15975
rect 16591 15941 16625 15975
rect 16659 15941 16693 15975
rect 16727 15941 16761 15975
rect 16795 15941 16829 15975
rect 16863 15941 16897 15975
rect 16931 15941 16965 15975
rect 16999 15941 17033 15975
rect 17067 15941 17101 15975
rect 17135 15941 17169 15975
rect 17239 15942 17273 15976
rect 17307 15942 17341 15976
rect 17375 15942 17409 15976
rect 17443 15942 17477 15976
rect 17511 15942 17545 15976
rect 17579 15942 17613 15976
rect 17647 15942 17681 15976
rect 17715 15942 17749 15976
rect 17783 15942 17817 15976
rect 17851 15942 17885 15976
rect 17919 15942 17953 15976
rect 17987 15942 18021 15976
rect 18055 15942 18089 15976
rect 15003 15868 15037 15902
rect 15003 15800 15037 15834
rect 15003 15732 15037 15766
rect 15003 15664 15037 15698
rect 15003 15596 15037 15630
rect 15003 15528 15037 15562
rect 15003 15460 15037 15494
rect 15003 15392 15037 15426
rect 15003 15324 15037 15358
rect 15003 15256 15037 15290
rect 15003 15188 15037 15222
rect 15003 15120 15037 15154
rect 15003 15052 15037 15086
rect 15003 14984 15037 15018
rect 15003 14916 15037 14950
rect 15003 14848 15037 14882
rect 18171 15918 18205 15952
rect 18171 15850 18205 15884
rect 18171 15782 18205 15816
rect 18171 15714 18205 15748
rect 18171 15646 18205 15680
rect 18171 15578 18205 15612
rect 18171 15510 18205 15544
rect 18171 15442 18205 15476
rect 18171 15374 18205 15408
rect 18171 15306 18205 15340
rect 18171 15238 18205 15272
rect 18171 15170 18205 15204
rect 18171 15102 18205 15136
rect 18171 15034 18205 15068
rect 18171 14966 18205 15000
rect 18171 14898 18205 14932
rect 15118 14824 15152 14858
rect 15186 14824 15220 14858
rect 15254 14824 15288 14858
rect 15322 14824 15356 14858
rect 15390 14824 15424 14858
rect 15458 14824 15492 14858
rect 15526 14824 15560 14858
rect 15594 14824 15628 14858
rect 15662 14824 15696 14858
rect 15730 14824 15764 14858
rect 15798 14824 15832 14858
rect 15866 14824 15900 14858
rect 15934 14824 15968 14858
rect 16002 14824 16036 14858
rect 16070 14824 16104 14858
rect 16138 14824 16172 14858
rect 16206 14824 16240 14858
rect 16274 14824 16308 14858
rect 16342 14824 16376 14858
rect 16410 14824 16444 14858
rect 16478 14824 16512 14858
rect 16546 14824 16580 14858
rect 16651 14824 16685 14858
rect 16719 14824 16753 14858
rect 16787 14824 16821 14858
rect 16855 14824 16889 14858
rect 16923 14824 16957 14858
rect 16991 14824 17025 14858
rect 17059 14824 17093 14858
rect 17127 14824 17161 14858
rect 17195 14824 17229 14858
rect 17263 14824 17297 14858
rect 17331 14824 17365 14858
rect 17399 14824 17433 14858
rect 17467 14824 17501 14858
rect 17535 14824 17569 14858
rect 17603 14824 17637 14858
rect 17671 14824 17705 14858
rect 17739 14824 17773 14858
rect 17807 14824 17841 14858
rect 17875 14824 17909 14858
rect 17943 14824 17977 14858
rect 18011 14824 18045 14858
rect 18079 14824 18113 14858
rect 18147 14824 18181 14858
<< poly >>
rect 9622 37386 10222 37416
rect 10384 37386 10984 37416
rect 11040 37386 11640 37416
rect 11696 37386 12296 37416
rect 12352 37386 12952 37416
rect 13008 37386 13608 37416
rect 13664 37386 14264 37416
rect 9622 35964 10222 36036
rect 10384 35964 10984 36036
rect 11040 35964 11640 36036
rect 11696 35964 12296 36036
rect 12352 35964 12952 36036
rect 13008 35964 13608 36036
rect 13664 35964 14264 36036
rect 14426 35984 15026 36017
rect 9622 34566 10222 34614
rect 9622 34532 9638 34566
rect 9672 34532 9714 34566
rect 9748 34532 9790 34566
rect 9824 34532 9866 34566
rect 9900 34532 9942 34566
rect 9976 34532 10018 34566
rect 10052 34532 10095 34566
rect 10129 34532 10172 34566
rect 10206 34532 10222 34566
rect 9622 34522 10222 34532
rect 10384 34566 10984 34614
rect 10384 34532 10400 34566
rect 10434 34532 10476 34566
rect 10510 34532 10552 34566
rect 10586 34532 10628 34566
rect 10662 34532 10704 34566
rect 10738 34532 10780 34566
rect 10814 34532 10857 34566
rect 10891 34532 10934 34566
rect 10968 34532 10984 34566
rect 10384 34522 10984 34532
rect 11040 34566 11640 34614
rect 11040 34532 11056 34566
rect 11090 34532 11132 34566
rect 11166 34532 11208 34566
rect 11242 34532 11284 34566
rect 11318 34532 11360 34566
rect 11394 34532 11436 34566
rect 11470 34532 11513 34566
rect 11547 34532 11590 34566
rect 11624 34532 11640 34566
rect 11040 34522 11640 34532
rect 11696 34566 12296 34614
rect 11696 34532 11712 34566
rect 11746 34532 11789 34566
rect 11823 34532 11866 34566
rect 11900 34532 11942 34566
rect 11976 34532 12018 34566
rect 12052 34532 12094 34566
rect 12128 34532 12170 34566
rect 12204 34532 12246 34566
rect 12280 34532 12296 34566
rect 11696 34522 12296 34532
rect 12352 34566 12952 34614
rect 12352 34532 12368 34566
rect 12402 34532 12444 34566
rect 12478 34532 12520 34566
rect 12554 34532 12596 34566
rect 12630 34532 12672 34566
rect 12706 34532 12748 34566
rect 12782 34532 12825 34566
rect 12859 34532 12902 34566
rect 12936 34532 12952 34566
rect 12352 34522 12952 34532
rect 13008 34566 13608 34614
rect 13008 34532 13024 34566
rect 13058 34532 13101 34566
rect 13135 34532 13178 34566
rect 13212 34532 13254 34566
rect 13288 34532 13330 34566
rect 13364 34532 13406 34566
rect 13440 34532 13482 34566
rect 13516 34532 13558 34566
rect 13592 34532 13608 34566
rect 13008 34522 13608 34532
rect 13664 34566 14264 34614
rect 13664 34532 13680 34566
rect 13714 34532 13757 34566
rect 13791 34532 13834 34566
rect 13868 34532 13910 34566
rect 13944 34532 13986 34566
rect 14020 34532 14062 34566
rect 14096 34532 14138 34566
rect 14172 34532 14214 34566
rect 14248 34532 14264 34566
rect 13664 34522 14264 34532
rect 19132 37368 19732 37398
rect 19788 37368 20388 37398
rect 20444 37368 21044 37398
rect 21100 37368 21700 37398
rect 21756 37368 22356 37398
rect 22412 37368 23012 37398
rect 19132 35988 19732 36018
rect 19788 35988 20388 36018
rect 20444 35988 21044 36018
rect 21100 35988 21700 36018
rect 21756 35988 22356 36018
rect 22412 35988 23012 36018
rect 9820 34181 10020 34191
rect 9820 34147 9836 34181
rect 9870 34147 9970 34181
rect 10004 34147 10020 34181
rect 9820 34099 10020 34147
rect 10076 34181 10276 34191
rect 10076 34147 10092 34181
rect 10126 34147 10226 34181
rect 10260 34147 10276 34181
rect 10076 34099 10276 34147
rect 10950 34181 11150 34191
rect 10950 34147 10966 34181
rect 11000 34147 11100 34181
rect 11134 34147 11150 34181
rect 10332 34099 10532 34129
rect 10694 34099 10894 34129
rect 10950 34099 11150 34147
rect 11206 34181 11406 34191
rect 11206 34147 11222 34181
rect 11256 34147 11356 34181
rect 11390 34147 11406 34181
rect 11206 34099 11406 34147
rect 8583 33644 8659 33663
rect 8280 33634 8430 33644
rect 8280 33600 8317 33634
rect 8351 33600 8430 33634
rect 8280 33584 8430 33600
rect 8583 33610 8606 33644
rect 8640 33610 8659 33644
rect 8583 33591 8659 33610
rect 8398 33476 8430 33584
rect 8607 33478 8637 33591
rect 8292 33446 8430 33476
rect 8606 33444 8738 33478
rect 9820 33451 10020 33499
rect 9820 33417 9836 33451
rect 9870 33417 9970 33451
rect 10004 33417 10020 33451
rect 9820 33407 10020 33417
rect 10076 33451 10276 33499
rect 10076 33417 10092 33451
rect 10126 33417 10226 33451
rect 10260 33417 10276 33451
rect 10076 33407 10276 33417
rect 10332 33451 10532 33499
rect 10332 33417 10348 33451
rect 10382 33417 10482 33451
rect 10516 33417 10532 33451
rect 10332 33407 10532 33417
rect 10694 33451 10894 33499
rect 10694 33417 10710 33451
rect 10744 33417 10844 33451
rect 10878 33417 10894 33451
rect 10694 33407 10894 33417
rect 10950 33451 11150 33499
rect 10950 33417 10966 33451
rect 11000 33417 11100 33451
rect 11134 33417 11150 33451
rect 10950 33407 11150 33417
rect 11206 33451 11406 33499
rect 11206 33417 11222 33451
rect 11256 33417 11356 33451
rect 11390 33417 11406 33451
rect 11206 33407 11406 33417
tri 8709 33213 8739 33214 sw
rect 8709 33200 8739 33213
rect 8060 33176 8136 33194
rect 8206 33176 8238 33194
rect 8293 33180 8323 33193
rect 8501 33186 8531 33199
rect 8060 33171 8238 33176
rect 8060 33137 8078 33171
rect 8112 33137 8238 33171
rect 8292 33152 8323 33180
rect 8060 33132 8238 33137
rect 8280 33136 8323 33152
rect 8426 33172 8531 33186
rect 8426 33138 8446 33172
rect 8480 33138 8531 33172
rect 8060 33116 8136 33132
rect 8207 33089 8237 33132
rect 8280 33112 8322 33136
rect 8426 33126 8531 33138
rect 8501 33121 8531 33126
rect 8694 33120 8739 33200
rect 8781 33121 8811 33193
rect 8988 33186 9018 33218
rect 12008 34124 12208 34154
rect 12264 34124 12464 34154
rect 12520 34124 12720 34154
rect 12008 33366 12208 33414
rect 12008 33332 12024 33366
rect 12058 33332 12158 33366
rect 12192 33332 12208 33366
rect 12008 33322 12208 33332
rect 12264 33366 12464 33414
rect 12264 33332 12280 33366
rect 12314 33332 12414 33366
rect 12448 33332 12464 33366
rect 12264 33322 12464 33332
rect 12520 33366 12720 33414
rect 12520 33332 12536 33366
rect 12570 33332 12670 33366
rect 12704 33332 12720 33366
rect 12520 33322 12720 33332
rect 19332 34258 19400 34324
rect 19351 34223 19381 34258
rect 13142 34106 13742 34136
rect 13920 34106 14520 34136
rect 19351 33902 19381 33963
rect 19330 33882 19400 33902
rect 19330 33848 19348 33882
rect 19382 33848 19400 33882
rect 19330 33830 19400 33848
rect 13142 33383 13742 33431
rect 13142 33349 13158 33383
rect 13192 33349 13234 33383
rect 13268 33349 13310 33383
rect 13344 33349 13386 33383
rect 13420 33349 13462 33383
rect 13496 33349 13538 33383
rect 13572 33349 13615 33383
rect 13649 33349 13692 33383
rect 13726 33349 13742 33383
rect 13142 33339 13742 33349
rect 13920 33383 14520 33431
rect 13920 33349 13936 33383
rect 13970 33349 14012 33383
rect 14046 33349 14088 33383
rect 14122 33349 14164 33383
rect 14198 33349 14240 33383
rect 14274 33349 14316 33383
rect 14350 33349 14393 33383
rect 14427 33349 14470 33383
rect 14504 33349 14520 33383
rect 13920 33339 14520 33349
rect 8906 33170 9018 33186
rect 8906 33136 8926 33170
rect 8960 33136 9018 33170
rect 8906 33126 9018 33136
rect 8988 33121 9018 33126
rect 7366 33002 7446 33024
rect 7366 32993 7903 33002
rect 7366 32959 7389 32993
rect 7423 32972 7903 32993
rect 7423 32959 7559 32972
rect 7366 32954 7559 32959
rect 7366 32934 7446 32954
rect 7529 32952 7559 32954
rect 7615 32950 7645 32972
rect 7701 32948 7731 32972
rect 7787 32932 7817 32972
rect 7873 32932 7903 32972
rect 8780 32844 8922 32874
rect 8886 32726 8922 32844
rect 9674 32794 9974 32824
rect 10030 32794 10330 32824
rect 10386 32794 10686 32824
rect 10742 32794 11042 32824
rect 8870 32710 8938 32726
rect 8870 32676 8886 32710
rect 8920 32676 8938 32710
rect 8870 32656 8938 32676
rect 11495 32930 11995 32940
rect 11495 32896 11511 32930
rect 11545 32896 11584 32930
rect 11618 32896 11657 32930
rect 11691 32896 11729 32930
rect 11763 32896 11801 32930
rect 11835 32896 11873 32930
rect 11907 32896 11945 32930
rect 11979 32896 11995 32930
rect 11495 32848 11995 32896
rect 12051 32930 12551 32940
rect 12051 32896 12067 32930
rect 12101 32896 12140 32930
rect 12174 32896 12213 32930
rect 12247 32896 12285 32930
rect 12319 32896 12357 32930
rect 12391 32896 12429 32930
rect 12463 32896 12501 32930
rect 12535 32896 12551 32930
rect 12051 32848 12551 32896
rect 12607 32930 13107 32940
rect 12607 32896 12623 32930
rect 12657 32896 12695 32930
rect 12729 32896 12767 32930
rect 12801 32896 12839 32930
rect 12873 32896 12911 32930
rect 12945 32896 12984 32930
rect 13018 32896 13057 32930
rect 13091 32896 13107 32930
rect 12607 32848 13107 32896
rect 13269 32930 13769 32940
rect 13269 32896 13285 32930
rect 13319 32896 13357 32930
rect 13391 32896 13429 32930
rect 13463 32896 13501 32930
rect 13535 32896 13573 32930
rect 13607 32896 13646 32930
rect 13680 32896 13719 32930
rect 13753 32896 13769 32930
rect 13269 32848 13769 32896
rect 13825 32930 14325 32940
rect 13825 32896 13841 32930
rect 13875 32896 13914 32930
rect 13948 32896 13987 32930
rect 14021 32896 14059 32930
rect 14093 32896 14131 32930
rect 14165 32896 14203 32930
rect 14237 32896 14275 32930
rect 14309 32896 14325 32930
rect 13825 32848 14325 32896
rect 11495 32294 11995 32348
rect 12051 32294 12551 32348
rect 12607 32294 13107 32348
rect 13269 32294 13769 32348
rect 13825 32294 14325 32348
rect 11495 31764 11995 31794
rect 12051 31764 12551 31794
rect 12607 31764 13107 31794
rect 13269 31764 13769 31794
rect 13825 31764 14325 31794
rect 9674 31346 9974 31394
rect 9674 31312 9690 31346
rect 9724 31312 9768 31346
rect 9802 31312 9846 31346
rect 9880 31312 9924 31346
rect 9958 31312 9974 31346
rect 9674 31302 9974 31312
rect 10030 31346 10330 31394
rect 10030 31312 10046 31346
rect 10080 31312 10124 31346
rect 10158 31312 10202 31346
rect 10236 31312 10280 31346
rect 10314 31312 10330 31346
rect 10030 31302 10330 31312
rect 10386 31346 10686 31394
rect 10386 31312 10402 31346
rect 10436 31312 10480 31346
rect 10514 31312 10558 31346
rect 10592 31312 10636 31346
rect 10670 31312 10686 31346
rect 10386 31302 10686 31312
rect 10742 31346 11042 31394
rect 10742 31312 10758 31346
rect 10792 31312 10836 31346
rect 10870 31312 10914 31346
rect 10948 31312 10992 31346
rect 11026 31312 11042 31346
rect 10742 31302 11042 31312
rect 9674 31162 9974 31172
rect 9674 31128 9690 31162
rect 9724 31128 9768 31162
rect 9802 31128 9846 31162
rect 9880 31128 9924 31162
rect 9958 31128 9974 31162
rect 9674 31080 9974 31128
rect 10030 31162 10330 31172
rect 10030 31128 10046 31162
rect 10080 31128 10124 31162
rect 10158 31128 10202 31162
rect 10236 31128 10280 31162
rect 10314 31128 10330 31162
rect 10030 31080 10330 31128
rect 10386 31162 10686 31172
rect 10386 31128 10402 31162
rect 10436 31128 10480 31162
rect 10514 31128 10558 31162
rect 10592 31128 10636 31162
rect 10670 31128 10686 31162
rect 10386 31080 10686 31128
rect 10742 31162 11042 31172
rect 10742 31128 10758 31162
rect 10792 31128 10836 31162
rect 10870 31128 10914 31162
rect 10948 31128 10992 31162
rect 11026 31128 11042 31162
rect 10742 31080 11042 31128
rect 11376 31190 11446 31206
rect 11376 31156 11396 31190
rect 11430 31188 11446 31190
rect 11430 31158 11492 31188
rect 11430 31156 11446 31158
rect 11376 31138 11446 31156
rect 9674 29650 9974 29680
rect 10030 29650 10330 29680
rect 10386 29650 10686 29680
rect 10742 29650 11042 29680
rect 11634 17608 12234 17641
rect 12396 17608 12996 17641
rect 13052 17608 13652 17641
rect 13708 17608 14308 17641
rect 14364 17608 14964 17641
rect 15020 17608 15620 17641
rect 15676 17608 16276 17641
rect 16438 17608 17038 17641
rect 10595 15268 10671 15287
rect 10292 15258 10442 15268
rect 10292 15224 10329 15258
rect 10363 15224 10442 15258
rect 10292 15208 10442 15224
rect 10595 15234 10618 15268
rect 10652 15234 10671 15268
rect 10595 15215 10671 15234
rect 10410 15100 10442 15208
rect 10619 15102 10649 15215
rect 10304 15070 10442 15100
rect 10618 15068 10750 15102
tri 10721 14837 10751 14838 sw
rect 10721 14824 10751 14837
rect 10072 14800 10148 14818
rect 10218 14800 10250 14818
rect 10305 14804 10335 14817
rect 10513 14810 10543 14823
rect 10072 14795 10250 14800
rect 10072 14761 10090 14795
rect 10124 14761 10250 14795
rect 10304 14776 10335 14804
rect 10072 14756 10250 14761
rect 10292 14760 10335 14776
rect 10438 14796 10543 14810
rect 10438 14762 10458 14796
rect 10492 14762 10543 14796
rect 10072 14740 10148 14756
rect 10219 14713 10249 14756
rect 10292 14736 10334 14760
rect 10438 14750 10543 14762
rect 10513 14745 10543 14750
rect 10706 14744 10751 14824
rect 10793 14745 10823 14817
rect 11000 14810 11030 14842
rect 21344 15882 21412 15948
rect 21363 15847 21393 15882
rect 21363 15526 21393 15587
rect 21342 15506 21412 15526
rect 21342 15472 21360 15506
rect 21394 15472 21412 15506
rect 21342 15454 21412 15472
rect 10918 14794 11030 14810
rect 10918 14760 10938 14794
rect 10972 14760 11030 14794
rect 10918 14750 11030 14760
rect 11000 14745 11030 14750
rect 9378 14626 9458 14648
rect 9378 14617 9915 14626
rect 9378 14583 9401 14617
rect 9435 14596 9915 14617
rect 9435 14583 9571 14596
rect 9378 14578 9571 14583
rect 9378 14558 9458 14578
rect 9541 14576 9571 14578
rect 9627 14574 9657 14596
rect 9713 14572 9743 14596
rect 9799 14556 9829 14596
rect 9885 14556 9915 14596
rect 10792 14468 10934 14498
rect 10898 14350 10934 14468
rect 10882 14334 10950 14350
rect 10882 14300 10898 14334
rect 10932 14300 10950 14334
rect 10882 14280 10950 14300
rect 13388 12814 13458 12830
rect 13388 12780 13408 12814
rect 13442 12812 13458 12814
rect 13442 12782 13504 12812
rect 13442 12780 13458 12782
rect 13388 12762 13458 12780
<< polycont >>
rect 9638 34532 9672 34566
rect 9714 34532 9748 34566
rect 9790 34532 9824 34566
rect 9866 34532 9900 34566
rect 9942 34532 9976 34566
rect 10018 34532 10052 34566
rect 10095 34532 10129 34566
rect 10172 34532 10206 34566
rect 10400 34532 10434 34566
rect 10476 34532 10510 34566
rect 10552 34532 10586 34566
rect 10628 34532 10662 34566
rect 10704 34532 10738 34566
rect 10780 34532 10814 34566
rect 10857 34532 10891 34566
rect 10934 34532 10968 34566
rect 11056 34532 11090 34566
rect 11132 34532 11166 34566
rect 11208 34532 11242 34566
rect 11284 34532 11318 34566
rect 11360 34532 11394 34566
rect 11436 34532 11470 34566
rect 11513 34532 11547 34566
rect 11590 34532 11624 34566
rect 11712 34532 11746 34566
rect 11789 34532 11823 34566
rect 11866 34532 11900 34566
rect 11942 34532 11976 34566
rect 12018 34532 12052 34566
rect 12094 34532 12128 34566
rect 12170 34532 12204 34566
rect 12246 34532 12280 34566
rect 12368 34532 12402 34566
rect 12444 34532 12478 34566
rect 12520 34532 12554 34566
rect 12596 34532 12630 34566
rect 12672 34532 12706 34566
rect 12748 34532 12782 34566
rect 12825 34532 12859 34566
rect 12902 34532 12936 34566
rect 13024 34532 13058 34566
rect 13101 34532 13135 34566
rect 13178 34532 13212 34566
rect 13254 34532 13288 34566
rect 13330 34532 13364 34566
rect 13406 34532 13440 34566
rect 13482 34532 13516 34566
rect 13558 34532 13592 34566
rect 13680 34532 13714 34566
rect 13757 34532 13791 34566
rect 13834 34532 13868 34566
rect 13910 34532 13944 34566
rect 13986 34532 14020 34566
rect 14062 34532 14096 34566
rect 14138 34532 14172 34566
rect 14214 34532 14248 34566
rect 9836 34147 9870 34181
rect 9970 34147 10004 34181
rect 10092 34147 10126 34181
rect 10226 34147 10260 34181
rect 10966 34147 11000 34181
rect 11100 34147 11134 34181
rect 11222 34147 11256 34181
rect 11356 34147 11390 34181
rect 8317 33600 8351 33634
rect 8606 33610 8640 33644
rect 9836 33417 9870 33451
rect 9970 33417 10004 33451
rect 10092 33417 10126 33451
rect 10226 33417 10260 33451
rect 10348 33417 10382 33451
rect 10482 33417 10516 33451
rect 10710 33417 10744 33451
rect 10844 33417 10878 33451
rect 10966 33417 11000 33451
rect 11100 33417 11134 33451
rect 11222 33417 11256 33451
rect 11356 33417 11390 33451
rect 8078 33137 8112 33171
rect 8446 33138 8480 33172
rect 12024 33332 12058 33366
rect 12158 33332 12192 33366
rect 12280 33332 12314 33366
rect 12414 33332 12448 33366
rect 12536 33332 12570 33366
rect 12670 33332 12704 33366
rect 19348 33848 19382 33882
rect 13158 33349 13192 33383
rect 13234 33349 13268 33383
rect 13310 33349 13344 33383
rect 13386 33349 13420 33383
rect 13462 33349 13496 33383
rect 13538 33349 13572 33383
rect 13615 33349 13649 33383
rect 13692 33349 13726 33383
rect 13936 33349 13970 33383
rect 14012 33349 14046 33383
rect 14088 33349 14122 33383
rect 14164 33349 14198 33383
rect 14240 33349 14274 33383
rect 14316 33349 14350 33383
rect 14393 33349 14427 33383
rect 14470 33349 14504 33383
rect 8926 33136 8960 33170
rect 7389 32959 7423 32993
rect 8886 32676 8920 32710
rect 11511 32896 11545 32930
rect 11584 32896 11618 32930
rect 11657 32896 11691 32930
rect 11729 32896 11763 32930
rect 11801 32896 11835 32930
rect 11873 32896 11907 32930
rect 11945 32896 11979 32930
rect 12067 32896 12101 32930
rect 12140 32896 12174 32930
rect 12213 32896 12247 32930
rect 12285 32896 12319 32930
rect 12357 32896 12391 32930
rect 12429 32896 12463 32930
rect 12501 32896 12535 32930
rect 12623 32896 12657 32930
rect 12695 32896 12729 32930
rect 12767 32896 12801 32930
rect 12839 32896 12873 32930
rect 12911 32896 12945 32930
rect 12984 32896 13018 32930
rect 13057 32896 13091 32930
rect 13285 32896 13319 32930
rect 13357 32896 13391 32930
rect 13429 32896 13463 32930
rect 13501 32896 13535 32930
rect 13573 32896 13607 32930
rect 13646 32896 13680 32930
rect 13719 32896 13753 32930
rect 13841 32896 13875 32930
rect 13914 32896 13948 32930
rect 13987 32896 14021 32930
rect 14059 32896 14093 32930
rect 14131 32896 14165 32930
rect 14203 32896 14237 32930
rect 14275 32896 14309 32930
rect 9690 31312 9724 31346
rect 9768 31312 9802 31346
rect 9846 31312 9880 31346
rect 9924 31312 9958 31346
rect 10046 31312 10080 31346
rect 10124 31312 10158 31346
rect 10202 31312 10236 31346
rect 10280 31312 10314 31346
rect 10402 31312 10436 31346
rect 10480 31312 10514 31346
rect 10558 31312 10592 31346
rect 10636 31312 10670 31346
rect 10758 31312 10792 31346
rect 10836 31312 10870 31346
rect 10914 31312 10948 31346
rect 10992 31312 11026 31346
rect 9690 31128 9724 31162
rect 9768 31128 9802 31162
rect 9846 31128 9880 31162
rect 9924 31128 9958 31162
rect 10046 31128 10080 31162
rect 10124 31128 10158 31162
rect 10202 31128 10236 31162
rect 10280 31128 10314 31162
rect 10402 31128 10436 31162
rect 10480 31128 10514 31162
rect 10558 31128 10592 31162
rect 10636 31128 10670 31162
rect 10758 31128 10792 31162
rect 10836 31128 10870 31162
rect 10914 31128 10948 31162
rect 10992 31128 11026 31162
rect 11396 31156 11430 31190
rect 10329 15224 10363 15258
rect 10618 15234 10652 15268
rect 10090 14761 10124 14795
rect 10458 14762 10492 14796
rect 21360 15472 21394 15506
rect 10938 14760 10972 14794
rect 9401 14583 9435 14617
rect 10898 14300 10932 14334
rect 13408 12780 13442 12814
<< xpolycontact >>
rect 21836 33376 22268 33658
rect 23356 33376 23788 33658
rect 21836 33046 22268 33328
rect 23356 33046 23788 33328
rect 21836 32716 22268 32998
rect 23356 32716 23788 32998
rect 21836 32384 22268 32666
rect 23356 32384 23788 32666
rect 21836 32056 22268 32338
rect 23356 32056 23788 32338
rect 21836 31726 22268 32008
rect 23356 31726 23788 32008
rect 21836 31396 22268 31678
rect 23356 31396 23788 31678
rect 12798 31180 13230 31250
rect 14058 31180 14490 31250
rect 21836 31066 22268 31348
rect 23356 31066 23788 31348
<< xpolyres >>
rect 22268 33376 23356 33658
rect 22268 33046 23356 33328
rect 22268 32716 23356 32998
rect 22268 32384 23356 32666
rect 22268 32056 23356 32338
rect 22268 31726 23356 32008
rect 22268 31396 23356 31678
rect 13230 31180 14058 31250
rect 22268 31066 23356 31348
<< locali >>
rect 9445 37602 9469 37636
rect 9503 37602 9537 37636
rect 9571 37602 9605 37636
rect 9639 37602 9673 37636
rect 9707 37602 9741 37636
rect 9775 37602 9809 37636
rect 9843 37602 9877 37636
rect 9911 37602 9945 37636
rect 9979 37602 10013 37636
rect 10047 37602 10081 37636
rect 10115 37602 10149 37636
rect 10183 37602 10217 37636
rect 10251 37602 10285 37636
rect 10319 37602 10353 37636
rect 10387 37602 10421 37636
rect 10455 37602 10489 37636
rect 10523 37602 10557 37636
rect 10591 37602 10625 37636
rect 10659 37602 10693 37636
rect 10727 37602 10761 37636
rect 10795 37602 10829 37636
rect 10863 37602 10897 37636
rect 10931 37602 10965 37636
rect 10999 37602 11033 37636
rect 11067 37602 11101 37636
rect 11135 37602 11169 37636
rect 11203 37602 11237 37636
rect 11271 37602 11305 37636
rect 11339 37602 11373 37636
rect 11407 37602 11441 37636
rect 11475 37602 11509 37636
rect 11543 37602 11577 37636
rect 11611 37602 11645 37636
rect 11679 37602 11713 37636
rect 11747 37602 11781 37636
rect 11815 37602 11849 37636
rect 11883 37602 11917 37636
rect 11951 37602 11985 37636
rect 12019 37602 12053 37636
rect 12087 37602 12121 37636
rect 12155 37602 12189 37636
rect 12223 37602 12257 37636
rect 12291 37602 12348 37636
rect 12382 37602 12416 37636
rect 12450 37602 12484 37636
rect 12518 37602 12552 37636
rect 12586 37602 12620 37636
rect 12654 37602 12688 37636
rect 12722 37602 12756 37636
rect 12790 37602 12824 37636
rect 12858 37602 12892 37636
rect 12926 37602 12960 37636
rect 12994 37602 13028 37636
rect 13062 37602 13096 37636
rect 13130 37602 13164 37636
rect 13198 37602 13232 37636
rect 13266 37602 13300 37636
rect 13334 37602 13368 37636
rect 13402 37602 13436 37636
rect 13470 37602 13504 37636
rect 13538 37602 13572 37636
rect 13606 37602 13640 37636
rect 13674 37602 13708 37636
rect 13742 37602 13776 37636
rect 13810 37602 13844 37636
rect 13878 37602 13912 37636
rect 13946 37602 13980 37636
rect 14014 37602 14048 37636
rect 14082 37602 14116 37636
rect 14150 37602 14184 37636
rect 14218 37602 14252 37636
rect 14286 37602 14320 37636
rect 14354 37602 14388 37636
rect 14422 37602 14456 37636
rect 14490 37602 14524 37636
rect 14558 37602 14592 37636
rect 14626 37602 14660 37636
rect 14694 37602 14728 37636
rect 14762 37602 14796 37636
rect 14830 37602 14864 37636
rect 14898 37602 14932 37636
rect 14966 37602 15000 37636
rect 15034 37602 15068 37636
rect 15102 37612 15371 37636
rect 15102 37602 15169 37612
rect 9445 37542 9479 37602
rect 15203 37578 15275 37612
rect 15309 37602 15371 37612
rect 15405 37602 15439 37636
rect 15473 37602 15507 37636
rect 15541 37602 15575 37636
rect 15609 37602 15643 37636
rect 15677 37602 15711 37636
rect 15745 37602 15779 37636
rect 15813 37602 15847 37636
rect 15881 37602 15915 37636
rect 15949 37602 15983 37636
rect 16017 37602 16051 37636
rect 16085 37602 16119 37636
rect 16153 37602 16187 37636
rect 16221 37602 16255 37636
rect 16289 37602 16323 37636
rect 16357 37602 16391 37636
rect 16425 37602 16459 37636
rect 16493 37602 16527 37636
rect 16561 37602 16595 37636
rect 16629 37602 16663 37636
rect 16697 37602 16731 37636
rect 16765 37602 16799 37636
rect 16833 37602 16867 37636
rect 16901 37602 16935 37636
rect 16969 37602 17003 37636
rect 17037 37602 17071 37636
rect 17105 37602 17139 37636
rect 17173 37602 17207 37636
rect 17241 37602 17275 37636
rect 17309 37602 17343 37636
rect 17377 37602 17411 37636
rect 17445 37602 17479 37636
rect 17513 37602 17547 37636
rect 17581 37602 17615 37636
rect 17649 37602 17683 37636
rect 17717 37602 17751 37636
rect 17785 37602 17819 37636
rect 17853 37602 17887 37636
rect 17921 37602 17955 37636
rect 17989 37602 18023 37636
rect 18057 37602 18091 37636
rect 18125 37602 18159 37636
rect 18193 37612 18362 37636
rect 18193 37602 18289 37612
rect 15169 37544 15309 37578
rect 15203 37510 15275 37544
rect 9479 37508 14401 37510
rect 9445 37500 14401 37508
rect 9445 37474 9599 37500
rect 9479 37466 9599 37474
rect 9651 37466 9667 37500
rect 9723 37466 9735 37500
rect 9795 37466 9803 37500
rect 9867 37466 9871 37500
rect 9973 37466 9977 37500
rect 10041 37466 10049 37500
rect 10109 37466 10121 37500
rect 10177 37466 10193 37500
rect 10245 37466 10358 37500
rect 10408 37466 10430 37500
rect 10476 37466 10502 37500
rect 10544 37466 10574 37500
rect 10612 37466 10646 37500
rect 10680 37466 10714 37500
rect 10752 37466 10782 37500
rect 10824 37466 10850 37500
rect 10896 37466 10918 37500
rect 10968 37466 11018 37500
rect 11068 37466 11090 37500
rect 11136 37466 11162 37500
rect 11204 37466 11234 37500
rect 11272 37466 11306 37500
rect 11340 37466 11374 37500
rect 11412 37466 11442 37500
rect 11484 37466 11510 37500
rect 11556 37466 11578 37500
rect 11628 37466 11674 37500
rect 11724 37466 11746 37500
rect 11792 37466 11818 37500
rect 11860 37466 11890 37500
rect 11928 37466 11962 37500
rect 11996 37466 12030 37500
rect 12068 37466 12098 37500
rect 12140 37466 12166 37500
rect 12212 37466 12234 37500
rect 12284 37466 12347 37500
rect 12397 37466 12419 37500
rect 12465 37466 12491 37500
rect 12533 37466 12563 37500
rect 12601 37466 12635 37500
rect 12669 37466 12703 37500
rect 12741 37466 12771 37500
rect 12813 37466 12839 37500
rect 12885 37466 12907 37500
rect 12957 37466 13020 37500
rect 13070 37466 13092 37500
rect 13138 37466 13164 37500
rect 13206 37466 13236 37500
rect 13274 37466 13308 37500
rect 13342 37466 13376 37500
rect 13414 37466 13444 37500
rect 13486 37466 13512 37500
rect 13558 37466 13580 37500
rect 13630 37466 13680 37500
rect 13730 37466 13752 37500
rect 13798 37466 13824 37500
rect 13866 37466 13896 37500
rect 13934 37466 13968 37500
rect 14002 37466 14036 37500
rect 14074 37466 14104 37500
rect 14146 37466 14172 37500
rect 14218 37466 14240 37500
rect 14290 37466 14401 37500
rect 9479 37456 14401 37466
rect 15072 37492 15309 37510
rect 18183 37578 18289 37602
rect 18323 37602 18362 37612
rect 18396 37602 18430 37636
rect 18464 37602 18498 37636
rect 18532 37602 18566 37636
rect 18600 37602 18634 37636
rect 18668 37602 18702 37636
rect 18736 37602 18770 37636
rect 18804 37602 18838 37636
rect 18872 37602 18906 37636
rect 18940 37602 18974 37636
rect 19008 37602 19042 37636
rect 19076 37602 19110 37636
rect 19144 37602 19178 37636
rect 19212 37602 19246 37636
rect 19280 37602 19314 37636
rect 19348 37602 19382 37636
rect 19416 37602 19450 37636
rect 19484 37602 19518 37636
rect 19552 37602 19586 37636
rect 19620 37602 19654 37636
rect 19688 37602 19722 37636
rect 19756 37602 19790 37636
rect 19824 37602 19858 37636
rect 19892 37602 19926 37636
rect 19960 37602 19994 37636
rect 20028 37602 20062 37636
rect 20096 37602 20130 37636
rect 20164 37602 20198 37636
rect 20232 37602 20266 37636
rect 20300 37602 20334 37636
rect 20368 37602 20402 37636
rect 20436 37602 20470 37636
rect 20504 37602 20538 37636
rect 20572 37602 20606 37636
rect 20640 37602 20674 37636
rect 20708 37602 20742 37636
rect 20776 37602 20810 37636
rect 20844 37602 20878 37636
rect 20912 37602 20946 37636
rect 20980 37602 21014 37636
rect 21048 37602 21145 37636
rect 21179 37602 21213 37636
rect 21247 37602 21281 37636
rect 21315 37602 21349 37636
rect 21383 37602 21417 37636
rect 21451 37602 21485 37636
rect 21519 37602 21553 37636
rect 21587 37602 21621 37636
rect 21655 37602 21689 37636
rect 21723 37602 21757 37636
rect 21791 37602 21825 37636
rect 21859 37602 21893 37636
rect 21927 37602 21961 37636
rect 21995 37602 22029 37636
rect 22063 37602 22097 37636
rect 22131 37602 22165 37636
rect 22199 37602 22233 37636
rect 22267 37602 22301 37636
rect 22335 37602 22369 37636
rect 22403 37602 22437 37636
rect 22471 37602 22505 37636
rect 22539 37602 22573 37636
rect 22607 37602 22641 37636
rect 22675 37602 22709 37636
rect 22743 37602 22777 37636
rect 22811 37602 22845 37636
rect 22879 37602 22913 37636
rect 22947 37602 22981 37636
rect 23015 37602 23049 37636
rect 23083 37602 23117 37636
rect 23151 37602 23185 37636
rect 23219 37602 23253 37636
rect 23287 37602 23321 37636
rect 23355 37602 23389 37636
rect 23423 37602 23457 37636
rect 23491 37602 23525 37636
rect 23559 37602 23593 37636
rect 23627 37602 23661 37636
rect 23695 37602 23729 37636
rect 23763 37602 23797 37636
rect 23831 37602 23855 37636
rect 18183 37544 18323 37578
rect 18183 37516 18289 37544
rect 15072 37476 15416 37492
rect 15072 37456 15169 37476
rect 9445 37406 9479 37440
rect 9445 37338 9479 37372
rect 9445 37270 9479 37304
rect 9445 37202 9479 37236
rect 9445 37134 9479 37168
rect 9445 37066 9479 37100
rect 9445 36998 9479 37032
rect 9445 36930 9479 36964
rect 9445 36862 9479 36896
rect 9445 36794 9479 36828
rect 9445 36726 9479 36760
rect 9445 36658 9479 36692
rect 9445 36590 9479 36624
rect 9445 36522 9479 36556
rect 9445 36454 9479 36488
rect 9445 36386 9479 36420
rect 9445 36318 9479 36352
rect 9445 36250 9479 36284
rect 9445 36182 9479 36216
rect 9445 36114 9479 36148
rect 9445 36046 9479 36080
rect 9445 35978 9479 36012
rect 9445 35910 9479 35944
rect 9445 35842 9479 35876
rect 9445 35774 9479 35808
rect 9445 35706 9479 35740
rect 9445 35638 9479 35672
rect 9445 35570 9479 35604
rect 9445 35502 9479 35536
rect 9445 35434 9479 35468
rect 9445 35366 9479 35400
rect 9445 35298 9479 35332
rect 9445 35230 9479 35264
rect 9445 35162 9479 35196
rect 9445 35094 9479 35128
rect 9445 35026 9479 35060
rect 9445 34958 9479 34992
rect 9445 34890 9479 34924
rect 9445 34822 9479 34856
rect 9445 34754 9479 34788
rect 6952 34688 6976 34722
rect 7010 34688 7044 34722
rect 7078 34688 7112 34722
rect 7146 34688 7180 34722
rect 7214 34688 7248 34722
rect 7282 34688 7316 34722
rect 7350 34688 7384 34722
rect 7418 34688 7452 34722
rect 7486 34688 7520 34722
rect 7554 34688 7588 34722
rect 7622 34688 7656 34722
rect 7690 34688 7724 34722
rect 7758 34688 7792 34722
rect 7826 34698 7926 34722
rect 7826 34688 7892 34698
rect 6952 34642 6986 34688
rect 6952 34574 6986 34608
rect 7892 34630 7926 34664
rect 7779 34596 7892 34597
rect 6952 34506 6986 34540
rect 6952 34438 6986 34472
rect 7452 34562 7926 34596
rect 7452 34528 7892 34562
rect 7452 34507 7926 34528
rect 7452 34506 7802 34507
rect 7452 34409 7562 34506
rect 7692 34409 7802 34506
rect 7892 34494 7926 34507
rect 7892 34426 7926 34460
rect 9445 34686 9479 34720
rect 9445 34618 9479 34652
rect 9577 37340 9611 37386
rect 9577 37272 9611 37306
rect 9577 37204 9611 37238
rect 9577 37136 9611 37170
rect 9577 37068 9611 37102
rect 9577 37000 9611 37034
rect 9577 36932 9611 36966
rect 9577 36864 9611 36898
rect 9577 36796 9611 36830
rect 9577 36728 9611 36762
rect 9577 36660 9611 36694
rect 9577 36592 9611 36626
rect 9577 36524 9611 36558
rect 9577 36456 9611 36490
rect 9577 36388 9611 36422
rect 9577 36320 9611 36354
rect 9577 36252 9611 36286
rect 9577 36184 9611 36218
rect 9577 36116 9611 36150
rect 9577 35918 9611 36082
rect 9577 35850 9611 35884
rect 9577 35782 9611 35816
rect 9577 35714 9611 35748
rect 9577 35646 9611 35680
rect 9577 35578 9611 35612
rect 9577 35510 9611 35544
rect 9577 35442 9611 35476
rect 9577 35374 9611 35408
rect 9577 35306 9611 35340
rect 9577 35238 9611 35272
rect 9577 35170 9611 35204
rect 9577 35102 9611 35136
rect 9577 35034 9611 35068
rect 9577 34966 9611 35000
rect 9577 34898 9611 34932
rect 9577 34830 9611 34864
rect 9577 34762 9611 34796
rect 9577 34694 9611 34728
rect 9577 34614 9611 34660
rect 10233 37340 10267 37386
rect 10233 37272 10267 37306
rect 10233 37204 10267 37238
rect 10233 37136 10267 37170
rect 10233 37068 10267 37102
rect 10233 37000 10267 37034
rect 10233 36932 10267 36966
rect 10233 36864 10267 36898
rect 10233 36796 10267 36830
rect 10233 36728 10267 36762
rect 10233 36660 10267 36694
rect 10233 36592 10267 36626
rect 10233 36524 10267 36558
rect 10233 36456 10267 36490
rect 10233 36388 10267 36422
rect 10233 36320 10267 36354
rect 10233 36252 10267 36286
rect 10233 36184 10267 36218
rect 10233 36116 10267 36150
rect 10233 35918 10267 36082
rect 10233 35850 10267 35884
rect 10233 35782 10267 35816
rect 10233 35714 10267 35748
rect 10233 35646 10267 35680
rect 10233 35578 10267 35612
rect 10233 35510 10267 35544
rect 10233 35442 10267 35476
rect 10233 35374 10267 35408
rect 10233 35306 10267 35340
rect 10233 35238 10267 35272
rect 10233 35170 10267 35204
rect 10233 35102 10267 35136
rect 10233 35034 10267 35068
rect 10233 34966 10267 35000
rect 10233 34898 10267 34932
rect 10233 34830 10267 34864
rect 10233 34762 10267 34796
rect 10233 34694 10267 34728
rect 10233 34614 10267 34660
rect 10339 37340 10373 37386
rect 10339 37272 10373 37306
rect 10339 37204 10373 37238
rect 10339 37136 10373 37170
rect 10339 37068 10373 37102
rect 10339 37000 10373 37034
rect 10339 36932 10373 36966
rect 10339 36864 10373 36898
rect 10339 36796 10373 36830
rect 10339 36728 10373 36762
rect 10339 36660 10373 36694
rect 10339 36592 10373 36626
rect 10339 36524 10373 36558
rect 10339 36456 10373 36490
rect 10339 36388 10373 36422
rect 10339 36320 10373 36354
rect 10339 36252 10373 36286
rect 10339 36184 10373 36218
rect 10339 36116 10373 36150
rect 10339 35918 10373 36082
rect 10339 35850 10373 35884
rect 10339 35782 10373 35816
rect 10339 35714 10373 35748
rect 10339 35646 10373 35680
rect 10339 35578 10373 35612
rect 10339 35510 10373 35544
rect 10339 35442 10373 35476
rect 10339 35374 10373 35408
rect 10339 35306 10373 35340
rect 10339 35238 10373 35272
rect 10339 35170 10373 35204
rect 10339 35102 10373 35136
rect 10339 35034 10373 35068
rect 10339 34966 10373 35000
rect 10339 34898 10373 34932
rect 10339 34830 10373 34864
rect 10339 34762 10373 34796
rect 10339 34694 10373 34728
rect 10339 34614 10373 34660
rect 10995 37340 11029 37386
rect 11650 37382 11686 37456
rect 10995 37272 11029 37306
rect 10995 37204 11029 37238
rect 10995 37136 11029 37170
rect 10995 37068 11029 37102
rect 10995 37000 11029 37034
rect 10995 36932 11029 36966
rect 10995 36864 11029 36898
rect 10995 36796 11029 36830
rect 10995 36728 11029 36762
rect 10995 36660 11029 36694
rect 10995 36592 11029 36626
rect 10995 36524 11029 36558
rect 10995 36456 11029 36490
rect 10995 36388 11029 36422
rect 10995 36320 11029 36354
rect 10995 36252 11029 36286
rect 10995 36184 11029 36218
rect 10995 36116 11029 36150
rect 10995 35918 11029 36082
rect 10995 35850 11029 35884
rect 10995 35782 11029 35816
rect 10995 35714 11029 35748
rect 10995 35646 11029 35680
rect 10995 35578 11029 35612
rect 10995 35510 11029 35544
rect 10995 35442 11029 35476
rect 10995 35374 11029 35408
rect 10995 35306 11029 35340
rect 10995 35238 11029 35272
rect 10995 35170 11029 35204
rect 10995 35102 11029 35136
rect 10995 35034 11029 35068
rect 10995 34966 11029 35000
rect 10995 34898 11029 34932
rect 10995 34830 11029 34864
rect 10995 34762 11029 34796
rect 10995 34694 11029 34728
rect 10995 34614 11029 34660
rect 11651 37340 11685 37382
rect 11651 37272 11685 37306
rect 11651 37204 11685 37238
rect 11651 37136 11685 37170
rect 11651 37068 11685 37102
rect 11651 37000 11685 37034
rect 11651 36932 11685 36966
rect 11651 36864 11685 36898
rect 11651 36796 11685 36830
rect 11651 36728 11685 36762
rect 11651 36660 11685 36694
rect 11651 36592 11685 36626
rect 11651 36524 11685 36558
rect 11651 36456 11685 36490
rect 11651 36388 11685 36422
rect 11651 36320 11685 36354
rect 11651 36252 11685 36286
rect 11651 36184 11685 36218
rect 11651 36116 11685 36150
rect 11651 35918 11685 36082
rect 11651 35850 11685 35884
rect 11651 35782 11685 35816
rect 11651 35714 11685 35748
rect 11651 35646 11685 35680
rect 11651 35578 11685 35612
rect 11651 35510 11685 35544
rect 11651 35442 11685 35476
rect 11651 35374 11685 35408
rect 11651 35306 11685 35340
rect 11651 35238 11685 35272
rect 11651 35170 11685 35204
rect 11651 35102 11685 35136
rect 11651 35034 11685 35068
rect 11651 34966 11685 35000
rect 11651 34898 11685 34932
rect 11651 34830 11685 34864
rect 11651 34762 11685 34796
rect 11651 34694 11685 34728
rect 11651 34614 11685 34660
rect 12307 37340 12341 37386
rect 12962 37380 12998 37456
rect 15203 37442 15275 37476
rect 15309 37442 15416 37476
rect 15169 37438 15416 37442
rect 16023 37438 16133 37492
rect 16691 37438 16801 37492
rect 17385 37438 17495 37492
rect 18077 37482 18183 37492
rect 18217 37510 18289 37516
rect 18217 37492 18323 37510
rect 23821 37542 23855 37602
rect 23821 37492 23855 37508
rect 18217 37482 18432 37492
rect 18077 37476 18432 37482
rect 18077 37448 18289 37476
rect 18077 37438 18183 37448
rect 15169 37408 15309 37438
rect 12307 37272 12341 37306
rect 12307 37204 12341 37238
rect 12307 37136 12341 37170
rect 12307 37068 12341 37102
rect 12307 37000 12341 37034
rect 12307 36932 12341 36966
rect 12307 36864 12341 36898
rect 12307 36796 12341 36830
rect 12307 36728 12341 36762
rect 12307 36660 12341 36694
rect 12307 36592 12341 36626
rect 12307 36524 12341 36558
rect 12307 36456 12341 36490
rect 12307 36388 12341 36422
rect 12307 36320 12341 36354
rect 12307 36252 12341 36286
rect 12307 36184 12341 36218
rect 12307 36116 12341 36150
rect 12307 35918 12341 36082
rect 12307 35850 12341 35884
rect 12307 35782 12341 35816
rect 12307 35714 12341 35748
rect 12307 35646 12341 35680
rect 12307 35578 12341 35612
rect 12307 35510 12341 35544
rect 12307 35442 12341 35476
rect 12307 35374 12341 35408
rect 12307 35306 12341 35340
rect 12307 35238 12341 35272
rect 12307 35170 12341 35204
rect 12307 35102 12341 35136
rect 12307 35034 12341 35068
rect 12307 34966 12341 35000
rect 12307 34898 12341 34932
rect 12307 34830 12341 34864
rect 12307 34762 12341 34796
rect 12307 34694 12341 34728
rect 12307 34614 12341 34660
rect 12963 37340 12997 37380
rect 12963 37272 12997 37306
rect 12963 37204 12997 37238
rect 12963 37136 12997 37170
rect 12963 37068 12997 37102
rect 12963 37000 12997 37034
rect 12963 36932 12997 36966
rect 12963 36864 12997 36898
rect 12963 36796 12997 36830
rect 12963 36728 12997 36762
rect 12963 36660 12997 36694
rect 12963 36592 12997 36626
rect 12963 36524 12997 36558
rect 12963 36456 12997 36490
rect 12963 36388 12997 36422
rect 12963 36320 12997 36354
rect 12963 36252 12997 36286
rect 12963 36184 12997 36218
rect 12963 36116 12997 36150
rect 12963 35918 12997 36082
rect 12963 35850 12997 35884
rect 12963 35782 12997 35816
rect 12963 35714 12997 35748
rect 12963 35646 12997 35680
rect 12963 35578 12997 35612
rect 12963 35510 12997 35544
rect 12963 35442 12997 35476
rect 12963 35374 12997 35408
rect 12963 35306 12997 35340
rect 12963 35238 12997 35272
rect 12963 35170 12997 35204
rect 12963 35102 12997 35136
rect 12963 35034 12997 35068
rect 12963 34966 12997 35000
rect 12963 34898 12997 34932
rect 12963 34830 12997 34864
rect 12963 34762 12997 34796
rect 12963 34694 12997 34728
rect 12963 34614 12997 34660
rect 13619 37340 13653 37386
rect 13619 37272 13653 37306
rect 13619 37204 13653 37238
rect 13619 37136 13653 37170
rect 13619 37068 13653 37102
rect 13619 37000 13653 37034
rect 13619 36932 13653 36966
rect 13619 36864 13653 36898
rect 13619 36796 13653 36830
rect 13619 36728 13653 36762
rect 13619 36660 13653 36694
rect 13619 36592 13653 36626
rect 13619 36524 13653 36558
rect 13619 36456 13653 36490
rect 13619 36388 13653 36422
rect 13619 36320 13653 36354
rect 13619 36252 13653 36286
rect 13619 36184 13653 36218
rect 13619 36116 13653 36150
rect 13619 35918 13653 36082
rect 13619 35850 13653 35884
rect 13619 35782 13653 35816
rect 13619 35714 13653 35748
rect 13619 35646 13653 35680
rect 13619 35578 13653 35612
rect 13619 35510 13653 35544
rect 13619 35442 13653 35476
rect 13619 35374 13653 35408
rect 13619 35306 13653 35340
rect 13619 35238 13653 35272
rect 13619 35170 13653 35204
rect 13619 35102 13653 35136
rect 13619 35034 13653 35068
rect 13619 34966 13653 35000
rect 13619 34898 13653 34932
rect 13619 34830 13653 34864
rect 13619 34762 13653 34796
rect 13619 34694 13653 34728
rect 13619 34614 13653 34660
rect 14275 37340 14309 37386
rect 14275 37272 14309 37306
rect 14275 37204 14309 37238
rect 14275 37136 14309 37170
rect 14275 37068 14309 37102
rect 14275 37000 14309 37034
rect 14275 36932 14309 36966
rect 14275 36864 14309 36898
rect 14275 36796 14309 36830
rect 14275 36728 14309 36762
rect 14275 36660 14309 36694
rect 14275 36592 14309 36626
rect 14275 36524 14309 36558
rect 14275 36456 14309 36490
rect 14275 36388 14309 36422
rect 14275 36320 14309 36354
rect 14275 36252 14309 36286
rect 14275 36184 14309 36218
rect 14275 36116 14309 36150
rect 14275 35918 14309 36082
rect 15203 37374 15275 37408
rect 15169 37340 15309 37374
rect 16728 37364 16764 37438
rect 18217 37442 18289 37448
rect 18323 37442 18432 37476
rect 18217 37438 18432 37442
rect 19042 37482 23131 37492
rect 19042 37448 19127 37482
rect 19177 37448 19199 37482
rect 19245 37448 19271 37482
rect 19313 37448 19343 37482
rect 19381 37448 19415 37482
rect 19449 37448 19483 37482
rect 19521 37448 19551 37482
rect 19593 37448 19619 37482
rect 19665 37448 19687 37482
rect 19737 37448 19800 37482
rect 19850 37448 19872 37482
rect 19918 37448 19944 37482
rect 19986 37448 20016 37482
rect 20054 37448 20088 37482
rect 20122 37448 20156 37482
rect 20194 37448 20224 37482
rect 20266 37448 20292 37482
rect 20338 37448 20360 37482
rect 20410 37448 20475 37482
rect 20523 37448 20547 37482
rect 20591 37448 20619 37482
rect 20659 37448 20691 37482
rect 20727 37448 20761 37482
rect 20797 37448 20829 37482
rect 20869 37448 20897 37482
rect 20941 37448 20965 37482
rect 21013 37448 21078 37482
rect 21128 37448 21150 37482
rect 21196 37448 21222 37482
rect 21264 37448 21294 37482
rect 21332 37448 21366 37482
rect 21400 37448 21434 37482
rect 21472 37448 21502 37482
rect 21544 37448 21570 37482
rect 21616 37448 21638 37482
rect 21688 37448 21751 37482
rect 21801 37448 21823 37482
rect 21869 37448 21895 37482
rect 21937 37448 21967 37482
rect 22005 37448 22039 37482
rect 22073 37448 22107 37482
rect 22145 37448 22175 37482
rect 22217 37448 22243 37482
rect 22289 37448 22311 37482
rect 22361 37448 22424 37482
rect 22474 37448 22496 37482
rect 22542 37448 22568 37482
rect 22610 37448 22640 37482
rect 22678 37448 22712 37482
rect 22746 37448 22780 37482
rect 22818 37448 22848 37482
rect 22890 37448 22916 37482
rect 22962 37448 22984 37482
rect 23034 37448 23131 37482
rect 19042 37438 23131 37448
rect 23715 37474 23855 37492
rect 23715 37440 23821 37474
rect 23715 37438 23855 37440
rect 18217 37414 18323 37438
rect 18183 37408 18323 37414
rect 18183 37380 18289 37408
rect 15203 37306 15275 37340
rect 15169 37272 15309 37306
rect 15203 37238 15275 37272
rect 15169 37204 15309 37238
rect 15203 37170 15275 37204
rect 15169 37136 15309 37170
rect 15203 37102 15275 37136
rect 15169 37068 15309 37102
rect 15203 37034 15275 37068
rect 15169 37000 15309 37034
rect 15203 36966 15275 37000
rect 15169 36932 15309 36966
rect 15203 36898 15275 36932
rect 15169 36864 15309 36898
rect 15203 36830 15275 36864
rect 15169 36796 15309 36830
rect 15203 36762 15275 36796
rect 15169 36728 15309 36762
rect 15203 36694 15275 36728
rect 15169 36660 15309 36694
rect 15203 36626 15275 36660
rect 15169 36592 15309 36626
rect 15203 36558 15275 36592
rect 15169 36524 15309 36558
rect 15203 36490 15275 36524
rect 15169 36456 15309 36490
rect 15203 36422 15275 36456
rect 15169 36388 15309 36422
rect 15203 36354 15275 36388
rect 15169 36320 15309 36354
rect 15203 36286 15275 36320
rect 15169 36252 15309 36286
rect 15203 36218 15275 36252
rect 15169 36184 15309 36218
rect 15203 36150 15275 36184
rect 15169 36116 15309 36150
rect 15203 36082 15275 36116
rect 18217 37374 18289 37380
rect 18217 37346 18323 37374
rect 18183 37340 18323 37346
rect 18183 37312 18289 37340
rect 18217 37306 18289 37312
rect 18217 37278 18323 37306
rect 18183 37272 18323 37278
rect 18183 37244 18289 37272
rect 18217 37238 18289 37244
rect 18217 37210 18323 37238
rect 18183 37204 18323 37210
rect 18183 37176 18289 37204
rect 18217 37170 18289 37176
rect 18217 37142 18323 37170
rect 18183 37136 18323 37142
rect 18183 37108 18289 37136
rect 18217 37102 18289 37108
rect 18217 37074 18323 37102
rect 18183 37068 18323 37074
rect 18183 37040 18289 37068
rect 18217 37034 18289 37040
rect 18217 37006 18323 37034
rect 18183 37000 18323 37006
rect 18183 36972 18289 37000
rect 18217 36966 18289 36972
rect 18217 36938 18323 36966
rect 18183 36932 18323 36938
rect 18183 36904 18289 36932
rect 18217 36898 18289 36904
rect 18217 36870 18323 36898
rect 18183 36864 18323 36870
rect 18183 36836 18289 36864
rect 18217 36830 18289 36836
rect 18217 36802 18323 36830
rect 18183 36796 18323 36802
rect 18183 36768 18289 36796
rect 18217 36762 18289 36768
rect 18217 36734 18323 36762
rect 18183 36728 18323 36734
rect 18183 36700 18289 36728
rect 18217 36694 18289 36700
rect 18217 36666 18323 36694
rect 18183 36660 18323 36666
rect 18183 36632 18289 36660
rect 18217 36626 18289 36632
rect 18217 36598 18323 36626
rect 18183 36592 18323 36598
rect 18183 36564 18289 36592
rect 18217 36558 18289 36564
rect 18217 36530 18323 36558
rect 18183 36524 18323 36530
rect 18183 36496 18289 36524
rect 18217 36490 18289 36496
rect 18217 36462 18323 36490
rect 18183 36456 18323 36462
rect 18183 36428 18289 36456
rect 18217 36422 18289 36428
rect 18217 36394 18323 36422
rect 18183 36388 18323 36394
rect 18183 36360 18289 36388
rect 18217 36354 18289 36360
rect 18217 36326 18323 36354
rect 18183 36320 18323 36326
rect 18183 36292 18289 36320
rect 18217 36286 18289 36292
rect 18217 36258 18323 36286
rect 18183 36252 18323 36258
rect 18183 36224 18289 36252
rect 18217 36218 18289 36224
rect 18217 36190 18323 36218
rect 18183 36184 18323 36190
rect 18183 36156 18289 36184
rect 18217 36150 18289 36156
rect 18217 36122 18323 36150
rect 18183 36116 18323 36122
rect 18183 36088 18289 36116
rect 15169 36048 15309 36082
rect 14381 35930 14415 36036
rect 15037 35930 15071 36036
rect 15203 36014 15275 36048
rect 15169 35980 15309 36014
rect 15203 35946 15275 35980
rect 14275 35850 14309 35884
rect 14275 35782 14309 35816
rect 14275 35714 14309 35748
rect 14275 35646 14309 35680
rect 14275 35578 14309 35612
rect 14275 35510 14309 35544
rect 14275 35442 14309 35476
rect 14275 35374 14309 35408
rect 14275 35306 14309 35340
rect 14275 35238 14309 35272
rect 14275 35170 14309 35204
rect 14275 35102 14309 35136
rect 14275 35034 14309 35068
rect 14275 34966 14309 35000
rect 14275 34898 14309 34932
rect 14275 34830 14309 34864
rect 14275 34762 14309 34796
rect 14275 34694 14309 34728
rect 14275 34614 14309 34660
rect 15169 35912 15309 35946
rect 15417 35930 15451 36018
rect 16073 35932 16107 36018
rect 16729 35930 16763 36084
rect 18217 36082 18289 36088
rect 18217 36054 18323 36082
rect 18183 36048 18323 36054
rect 19087 37322 19121 37368
rect 19087 37254 19121 37288
rect 19087 37186 19121 37220
rect 19087 37118 19121 37152
rect 19087 37050 19121 37084
rect 19087 36982 19121 37016
rect 19087 36914 19121 36948
rect 19087 36846 19121 36880
rect 19087 36778 19121 36812
rect 19087 36710 19121 36744
rect 19087 36642 19121 36676
rect 19087 36574 19121 36608
rect 19087 36506 19121 36540
rect 19087 36438 19121 36472
rect 19087 36370 19121 36404
rect 19087 36302 19121 36336
rect 19087 36234 19121 36268
rect 19087 36166 19121 36200
rect 19087 36098 19121 36132
rect 17385 35930 17419 36027
rect 18041 35930 18075 36027
rect 18183 36014 18289 36048
rect 18183 35980 18323 36014
rect 18183 35978 18289 35980
rect 18217 35946 18289 35978
rect 18431 35964 18465 36052
rect 19087 35964 19121 36064
rect 19743 37322 19777 37438
rect 19743 37254 19777 37288
rect 19743 37186 19777 37220
rect 19743 37118 19777 37152
rect 19743 37050 19777 37084
rect 19743 36982 19777 37016
rect 19743 36914 19777 36948
rect 19743 36846 19777 36880
rect 19743 36778 19777 36812
rect 19743 36710 19777 36744
rect 19743 36642 19777 36676
rect 19743 36574 19777 36608
rect 19743 36506 19777 36540
rect 19743 36438 19777 36472
rect 19743 36370 19777 36404
rect 19743 36302 19777 36336
rect 19743 36234 19777 36268
rect 19743 36166 19777 36200
rect 19743 36098 19777 36132
rect 19743 35964 19777 36064
rect 20399 37322 20433 37368
rect 20399 37254 20433 37288
rect 20399 37186 20433 37220
rect 20399 37118 20433 37152
rect 20399 37050 20433 37084
rect 20399 36982 20433 37016
rect 20399 36914 20433 36948
rect 20399 36846 20433 36880
rect 20399 36778 20433 36812
rect 20399 36710 20433 36744
rect 20399 36642 20433 36676
rect 20399 36574 20433 36608
rect 20399 36506 20433 36540
rect 20399 36438 20433 36472
rect 20399 36370 20433 36404
rect 20399 36302 20433 36336
rect 20399 36234 20433 36268
rect 20399 36166 20433 36200
rect 20399 36098 20433 36132
rect 20399 35964 20433 36064
rect 21055 37322 21089 37368
rect 21710 37358 21746 37438
rect 21055 37254 21089 37288
rect 21055 37186 21089 37220
rect 21055 37118 21089 37152
rect 21055 37050 21089 37084
rect 21055 36982 21089 37016
rect 21055 36914 21089 36948
rect 21055 36846 21089 36880
rect 21055 36778 21089 36812
rect 21055 36710 21089 36744
rect 21055 36642 21089 36676
rect 21055 36574 21089 36608
rect 21055 36506 21089 36540
rect 21055 36438 21089 36472
rect 21055 36370 21089 36404
rect 21055 36302 21089 36336
rect 21055 36234 21089 36268
rect 21055 36166 21089 36200
rect 21055 36098 21089 36132
rect 21055 35964 21089 36064
rect 21711 37322 21745 37358
rect 21711 37254 21745 37288
rect 21711 37186 21745 37220
rect 21711 37118 21745 37152
rect 21711 37050 21745 37084
rect 21711 36982 21745 37016
rect 21711 36914 21745 36948
rect 21711 36846 21745 36880
rect 21711 36778 21745 36812
rect 21711 36710 21745 36744
rect 21711 36642 21745 36676
rect 21711 36574 21745 36608
rect 21711 36506 21745 36540
rect 21711 36438 21745 36472
rect 21711 36370 21745 36404
rect 21711 36302 21745 36336
rect 21711 36234 21745 36268
rect 21711 36166 21745 36200
rect 21711 36098 21745 36132
rect 21711 35964 21745 36064
rect 22367 37322 22401 37368
rect 23022 37354 23058 37438
rect 23821 37406 23855 37438
rect 22367 37254 22401 37288
rect 22367 37186 22401 37220
rect 22367 37118 22401 37152
rect 22367 37050 22401 37084
rect 22367 36982 22401 37016
rect 22367 36914 22401 36948
rect 22367 36846 22401 36880
rect 22367 36778 22401 36812
rect 22367 36710 22401 36744
rect 22367 36642 22401 36676
rect 22367 36574 22401 36608
rect 22367 36506 22401 36540
rect 22367 36438 22401 36472
rect 22367 36370 22401 36404
rect 22367 36302 22401 36336
rect 22367 36234 22401 36268
rect 22367 36166 22401 36200
rect 22367 36098 22401 36132
rect 22367 35964 22401 36064
rect 23023 37322 23057 37354
rect 23023 37254 23057 37288
rect 23023 37186 23057 37220
rect 23023 37118 23057 37152
rect 23023 37050 23057 37084
rect 23023 36982 23057 37016
rect 23023 36914 23057 36948
rect 23023 36846 23057 36880
rect 23023 36778 23057 36812
rect 23023 36710 23057 36744
rect 23023 36642 23057 36676
rect 23023 36574 23057 36608
rect 23023 36506 23057 36540
rect 23023 36438 23057 36472
rect 23023 36370 23057 36404
rect 23023 36302 23057 36336
rect 23023 36234 23057 36268
rect 23023 36166 23057 36200
rect 23023 36098 23057 36132
rect 23023 35964 23057 36064
rect 23821 37338 23855 37372
rect 23821 37270 23855 37304
rect 23821 37202 23855 37236
rect 23821 37134 23855 37168
rect 23821 37066 23855 37100
rect 23821 36998 23855 37032
rect 23821 36930 23855 36964
rect 23821 36862 23855 36896
rect 23821 36794 23855 36828
rect 23821 36726 23855 36760
rect 23821 36658 23855 36692
rect 23821 36590 23855 36624
rect 23821 36522 23855 36556
rect 23821 36454 23855 36488
rect 23821 36386 23855 36420
rect 23821 36318 23855 36352
rect 23821 36250 23855 36284
rect 23821 36182 23855 36216
rect 23821 36114 23855 36148
rect 23679 35964 23713 36050
rect 23821 36046 23855 36080
rect 23821 35978 23855 36012
rect 18217 35944 18323 35946
rect 15203 35878 15275 35912
rect 15169 35844 15309 35878
rect 15203 35810 15275 35844
rect 15169 35776 15309 35810
rect 15203 35742 15275 35776
rect 15169 35708 15309 35742
rect 15203 35674 15275 35708
rect 15169 35640 15309 35674
rect 15203 35606 15275 35640
rect 15169 35572 15309 35606
rect 15203 35538 15275 35572
rect 15169 35504 15309 35538
rect 15203 35470 15275 35504
rect 15169 35436 15309 35470
rect 15203 35402 15275 35436
rect 15169 35368 15309 35402
rect 15203 35334 15275 35368
rect 15169 35300 15309 35334
rect 15203 35266 15275 35300
rect 15169 35232 15309 35266
rect 15203 35198 15275 35232
rect 15169 35164 15309 35198
rect 15203 35130 15275 35164
rect 15169 35096 15309 35130
rect 15203 35062 15275 35096
rect 15169 35028 15309 35062
rect 15203 34994 15275 35028
rect 15169 34960 15309 34994
rect 15203 34926 15275 34960
rect 15169 34892 15309 34926
rect 15203 34858 15275 34892
rect 18183 35912 18323 35944
rect 18183 35910 18289 35912
rect 18217 35878 18289 35910
rect 18217 35876 18323 35878
rect 18183 35844 18323 35876
rect 18183 35842 18289 35844
rect 18217 35810 18289 35842
rect 18217 35808 18323 35810
rect 18183 35776 18323 35808
rect 18183 35774 18289 35776
rect 18217 35742 18289 35774
rect 18217 35740 18323 35742
rect 18183 35708 18323 35740
rect 18183 35706 18289 35708
rect 18217 35674 18289 35706
rect 18217 35672 18323 35674
rect 18183 35640 18323 35672
rect 18183 35638 18289 35640
rect 18217 35606 18289 35638
rect 18217 35604 18323 35606
rect 18183 35572 18323 35604
rect 18183 35570 18289 35572
rect 18217 35538 18289 35570
rect 18217 35536 18323 35538
rect 18183 35504 18323 35536
rect 18183 35502 18289 35504
rect 18217 35470 18289 35502
rect 18217 35468 18323 35470
rect 18183 35436 18323 35468
rect 18183 35434 18289 35436
rect 18217 35402 18289 35434
rect 18217 35400 18323 35402
rect 18183 35368 18323 35400
rect 18183 35366 18289 35368
rect 18217 35334 18289 35366
rect 18217 35332 18323 35334
rect 18183 35300 18323 35332
rect 18183 35298 18289 35300
rect 18217 35266 18289 35298
rect 18217 35264 18323 35266
rect 18183 35232 18323 35264
rect 18183 35230 18289 35232
rect 18217 35198 18289 35230
rect 18217 35196 18323 35198
rect 18183 35164 18323 35196
rect 18183 35162 18289 35164
rect 18217 35130 18289 35162
rect 23821 35910 23855 35944
rect 23821 35842 23855 35876
rect 23821 35774 23855 35808
rect 23821 35706 23855 35740
rect 23821 35638 23855 35672
rect 23821 35570 23855 35604
rect 23821 35502 23855 35536
rect 23821 35434 23855 35468
rect 23821 35366 23855 35400
rect 23821 35298 23855 35332
rect 23821 35230 23855 35264
rect 23821 35162 23855 35196
rect 18217 35128 18323 35130
rect 18183 35096 18323 35128
rect 18183 35094 18289 35096
rect 18217 35062 18289 35094
rect 18217 35060 18323 35062
rect 18183 35028 18323 35060
rect 18183 35026 18289 35028
rect 18217 34994 18289 35026
rect 18217 34992 18323 34994
rect 18183 34960 18323 34992
rect 23679 34961 23713 35144
rect 23821 35094 23855 35128
rect 23821 35026 23855 35060
rect 18183 34958 18289 34960
rect 18217 34926 18289 34958
rect 18217 34924 18323 34926
rect 18183 34892 18323 34924
rect 18183 34890 18289 34892
rect 15169 34824 15309 34858
rect 15203 34790 15275 34824
rect 15169 34756 15309 34790
rect 15203 34722 15275 34756
rect 15169 34688 15309 34722
rect 15203 34654 15275 34688
rect 18041 34669 18075 34880
rect 18217 34858 18289 34890
rect 18217 34856 18323 34858
rect 18183 34824 18323 34856
rect 18183 34822 18289 34824
rect 18217 34790 18289 34822
rect 18217 34788 18323 34790
rect 18183 34756 18323 34788
rect 18183 34754 18289 34756
rect 18217 34722 18289 34754
rect 18217 34720 18323 34722
rect 18183 34688 18323 34720
rect 18183 34686 18289 34688
rect 15169 34620 15309 34654
rect 9445 34550 9479 34584
rect 15203 34586 15275 34620
rect 9622 34566 10222 34572
rect 9622 34532 9638 34566
rect 9672 34532 9714 34566
rect 9748 34532 9790 34566
rect 9824 34532 9866 34566
rect 9900 34532 9942 34566
rect 9976 34532 10018 34566
rect 10052 34532 10095 34566
rect 10129 34532 10172 34566
rect 10206 34532 10222 34566
rect 9622 34526 10222 34532
rect 10384 34566 10984 34572
rect 10384 34532 10400 34566
rect 10434 34532 10476 34566
rect 10510 34532 10552 34566
rect 10586 34532 10628 34566
rect 10662 34532 10704 34566
rect 10738 34532 10780 34566
rect 10814 34532 10857 34566
rect 10891 34532 10934 34566
rect 10968 34532 10984 34566
rect 10384 34526 10984 34532
rect 11040 34566 11640 34572
rect 11040 34532 11056 34566
rect 11090 34532 11132 34566
rect 11166 34532 11208 34566
rect 11242 34532 11284 34566
rect 11318 34532 11360 34566
rect 11394 34532 11436 34566
rect 11470 34532 11513 34566
rect 11547 34532 11590 34566
rect 11624 34532 11640 34566
rect 11040 34526 11640 34532
rect 11696 34566 12296 34572
rect 11696 34532 11712 34566
rect 11746 34532 11789 34566
rect 11823 34532 11866 34566
rect 11900 34532 11942 34566
rect 11976 34532 12018 34566
rect 12052 34532 12094 34566
rect 12128 34532 12170 34566
rect 12204 34532 12246 34566
rect 12280 34532 12296 34566
rect 11696 34526 12296 34532
rect 12352 34566 12952 34572
rect 12352 34532 12368 34566
rect 12402 34532 12444 34566
rect 12478 34532 12520 34566
rect 12554 34532 12596 34566
rect 12630 34532 12672 34566
rect 12706 34532 12748 34566
rect 12782 34532 12825 34566
rect 12859 34532 12902 34566
rect 12936 34532 12952 34566
rect 12352 34526 12952 34532
rect 13008 34566 13608 34572
rect 13008 34532 13024 34566
rect 13058 34532 13101 34566
rect 13135 34532 13178 34566
rect 13212 34532 13254 34566
rect 13288 34532 13330 34566
rect 13364 34532 13406 34566
rect 13440 34532 13482 34566
rect 13516 34532 13558 34566
rect 13592 34532 13608 34566
rect 13008 34526 13608 34532
rect 13664 34566 14264 34572
rect 13664 34532 13680 34566
rect 13714 34532 13757 34566
rect 13791 34532 13834 34566
rect 13868 34532 13910 34566
rect 13944 34532 13986 34566
rect 14020 34532 14062 34566
rect 14096 34532 14138 34566
rect 14172 34532 14214 34566
rect 14248 34532 14264 34566
rect 13664 34526 14264 34532
rect 15169 34552 15309 34586
rect 9445 34482 9479 34516
rect 15203 34518 15275 34552
rect 15169 34458 15309 34518
rect 18217 34654 18289 34686
rect 18217 34652 18323 34654
rect 18183 34620 18323 34652
rect 18183 34618 18289 34620
rect 18217 34586 18289 34618
rect 23821 34958 23855 34992
rect 23821 34890 23855 34924
rect 23821 34822 23855 34856
rect 23821 34754 23855 34788
rect 23821 34686 23855 34720
rect 23821 34618 23855 34652
rect 18217 34584 18323 34586
rect 18183 34552 18323 34584
rect 22367 34572 22401 34614
rect 18183 34550 18289 34552
rect 18217 34518 18289 34550
rect 22356 34526 22412 34572
rect 23821 34550 23855 34584
rect 18217 34516 18323 34518
rect 18183 34482 18323 34516
rect 9479 34448 9569 34458
rect 9445 34440 9569 34448
rect 6952 34370 6986 34404
rect 6952 34302 6986 34336
rect 6952 34234 6986 34268
rect 6952 34166 6986 34200
rect 6952 34098 6986 34132
rect 6952 34030 6986 34064
rect 6952 33891 6986 33996
rect 6952 33823 6986 33857
rect 6952 33755 6986 33789
rect 6952 33687 6986 33721
rect 6952 33619 6986 33653
rect 7892 34358 7926 34392
rect 7892 34290 7926 34324
rect 9266 34424 9569 34440
rect 9603 34424 9637 34458
rect 9671 34424 9705 34458
rect 9739 34424 9773 34458
rect 9807 34424 9841 34458
rect 9875 34424 9909 34458
rect 9943 34424 9977 34458
rect 10011 34424 10045 34458
rect 10079 34424 10113 34458
rect 10147 34424 10181 34458
rect 10215 34424 10249 34458
rect 10283 34424 10317 34458
rect 10351 34424 10385 34458
rect 10419 34424 10453 34458
rect 10487 34424 10521 34458
rect 10555 34424 10589 34458
rect 10623 34424 10657 34458
rect 10691 34424 10725 34458
rect 10759 34424 10793 34458
rect 10827 34424 10861 34458
rect 10895 34424 10929 34458
rect 10963 34424 10997 34458
rect 11031 34424 11065 34458
rect 11099 34424 11133 34458
rect 11167 34424 11201 34458
rect 11235 34424 11269 34458
rect 11303 34424 11337 34458
rect 11371 34424 11405 34458
rect 11439 34424 11473 34458
rect 11507 34424 11541 34458
rect 11575 34424 11609 34458
rect 11643 34424 11677 34458
rect 11711 34424 11745 34458
rect 11779 34424 11813 34458
rect 11847 34424 11881 34458
rect 11915 34424 11949 34458
rect 11983 34424 12017 34458
rect 12051 34424 12085 34458
rect 12119 34424 12153 34458
rect 12187 34424 12221 34458
rect 12255 34424 12289 34458
rect 12323 34424 12357 34458
rect 12391 34424 12425 34458
rect 12459 34424 12493 34458
rect 12527 34424 12561 34458
rect 12595 34424 12629 34458
rect 12663 34424 12697 34458
rect 12731 34424 12765 34458
rect 12799 34424 12833 34458
rect 12867 34424 12901 34458
rect 12935 34424 12969 34458
rect 13003 34424 13037 34458
rect 13071 34424 13105 34458
rect 13139 34424 13173 34458
rect 13207 34424 13241 34458
rect 13275 34424 13309 34458
rect 13343 34424 13377 34458
rect 13411 34424 13445 34458
rect 13479 34424 13513 34458
rect 13547 34424 13581 34458
rect 13615 34424 13649 34458
rect 13683 34424 13717 34458
rect 13751 34424 13785 34458
rect 13819 34424 13853 34458
rect 13887 34424 13921 34458
rect 13955 34424 13989 34458
rect 14023 34424 14057 34458
rect 14091 34424 14125 34458
rect 14159 34424 14193 34458
rect 14227 34424 14261 34458
rect 14295 34424 14329 34458
rect 14363 34424 14397 34458
rect 14431 34424 14465 34458
rect 14499 34424 14533 34458
rect 14567 34424 14601 34458
rect 14635 34424 14669 34458
rect 14703 34424 14737 34458
rect 14771 34424 14805 34458
rect 14839 34424 14873 34458
rect 14907 34424 14941 34458
rect 14975 34424 15009 34458
rect 15043 34424 15077 34458
rect 15111 34424 15145 34458
rect 15179 34424 15299 34458
rect 15333 34424 15367 34458
rect 15401 34424 15435 34458
rect 15469 34424 15503 34458
rect 15537 34424 15571 34458
rect 15605 34424 15639 34458
rect 15673 34424 15707 34458
rect 15741 34424 15775 34458
rect 15809 34424 15843 34458
rect 15877 34424 15911 34458
rect 15945 34424 15979 34458
rect 16013 34424 16047 34458
rect 16081 34424 16115 34458
rect 16149 34424 16183 34458
rect 16217 34424 16251 34458
rect 16285 34424 16319 34458
rect 16353 34424 16387 34458
rect 16421 34424 16455 34458
rect 16489 34424 16523 34458
rect 16557 34424 16591 34458
rect 16625 34424 16659 34458
rect 16693 34424 16727 34458
rect 16761 34424 16795 34458
rect 16829 34424 16863 34458
rect 16897 34424 16931 34458
rect 16965 34424 16999 34458
rect 17033 34424 17067 34458
rect 17101 34424 17135 34458
rect 17169 34424 17203 34458
rect 17237 34424 17271 34458
rect 17305 34424 17339 34458
rect 17373 34424 17407 34458
rect 17441 34424 17475 34458
rect 17509 34424 17543 34458
rect 17577 34424 17611 34458
rect 17645 34424 17679 34458
rect 17713 34424 17747 34458
rect 17781 34424 17815 34458
rect 17849 34424 17883 34458
rect 17917 34424 17951 34458
rect 17985 34424 18019 34458
rect 18053 34424 18087 34458
rect 18121 34448 18183 34458
rect 18217 34458 18323 34482
rect 23821 34482 23855 34516
rect 18217 34448 18313 34458
rect 18121 34424 18313 34448
rect 18347 34424 18381 34458
rect 18415 34424 18449 34458
rect 18483 34424 18517 34458
rect 18551 34424 18585 34458
rect 18619 34424 18653 34458
rect 18687 34424 18721 34458
rect 18755 34424 18789 34458
rect 18823 34424 18857 34458
rect 18891 34424 18925 34458
rect 18959 34424 18993 34458
rect 19027 34424 19061 34458
rect 19095 34424 19129 34458
rect 19163 34424 19197 34458
rect 19231 34424 19265 34458
rect 19299 34424 19333 34458
rect 19367 34424 19401 34458
rect 19435 34424 19469 34458
rect 19503 34424 19537 34458
rect 19571 34424 19605 34458
rect 19639 34424 19673 34458
rect 19707 34424 19741 34458
rect 19775 34424 19809 34458
rect 19843 34424 19877 34458
rect 19911 34424 19945 34458
rect 19979 34424 20013 34458
rect 20047 34424 20081 34458
rect 20115 34424 20149 34458
rect 20183 34424 20217 34458
rect 20251 34424 20285 34458
rect 20319 34424 20353 34458
rect 20387 34424 20421 34458
rect 20455 34424 20489 34458
rect 20523 34424 20557 34458
rect 20591 34424 20625 34458
rect 20659 34424 20693 34458
rect 20727 34424 20761 34458
rect 20795 34424 20829 34458
rect 20863 34424 20897 34458
rect 20931 34424 20965 34458
rect 20999 34424 21033 34458
rect 21067 34424 21101 34458
rect 21135 34424 21169 34458
rect 21203 34424 21237 34458
rect 21271 34424 21305 34458
rect 21339 34424 21373 34458
rect 21407 34424 21441 34458
rect 21475 34424 21509 34458
rect 21543 34424 21577 34458
rect 21611 34424 21645 34458
rect 21679 34424 21713 34458
rect 21747 34424 21781 34458
rect 21815 34424 21849 34458
rect 21883 34424 21917 34458
rect 21951 34424 21985 34458
rect 22019 34424 22053 34458
rect 22087 34424 22121 34458
rect 22155 34424 22189 34458
rect 22223 34424 22257 34458
rect 22291 34424 22325 34458
rect 22359 34424 22393 34458
rect 22427 34424 22461 34458
rect 22495 34424 22529 34458
rect 22563 34424 22597 34458
rect 22631 34424 22665 34458
rect 22699 34424 22733 34458
rect 22767 34424 22801 34458
rect 22835 34424 22869 34458
rect 22903 34424 22937 34458
rect 22971 34424 23005 34458
rect 23039 34424 23073 34458
rect 23107 34424 23141 34458
rect 23175 34424 23209 34458
rect 23243 34424 23277 34458
rect 23311 34424 23345 34458
rect 23379 34424 23413 34458
rect 23447 34424 23481 34458
rect 23515 34424 23549 34458
rect 23583 34424 23617 34458
rect 23651 34424 23685 34458
rect 23719 34424 23753 34458
rect 23787 34448 23821 34458
rect 23787 34424 23855 34448
rect 9266 34398 9504 34424
rect 9266 34364 9289 34398
rect 9323 34364 9504 34398
rect 9266 34352 9504 34364
rect 11692 34352 11750 34424
rect 9266 34322 9469 34352
rect 7892 34222 7926 34256
rect 7892 34154 7926 34188
rect 7892 34086 7926 34120
rect 7892 34018 7926 34052
rect 7892 33950 7926 33984
rect 7892 33882 7926 33916
rect 7892 33814 7926 33848
rect 7892 33746 7926 33780
rect 7892 33678 7926 33712
rect 9445 34318 9469 34322
rect 9503 34318 9537 34352
rect 9571 34318 9605 34352
rect 9639 34318 9673 34352
rect 9707 34318 9741 34352
rect 9775 34318 9809 34352
rect 9843 34318 9877 34352
rect 9911 34318 9945 34352
rect 9979 34318 10013 34352
rect 10047 34318 10081 34352
rect 10115 34318 10149 34352
rect 10183 34318 10217 34352
rect 10251 34318 10285 34352
rect 10319 34318 10353 34352
rect 10387 34318 10421 34352
rect 10455 34318 10489 34352
rect 10523 34318 10637 34352
rect 10671 34318 10705 34352
rect 10739 34318 10773 34352
rect 10807 34318 10841 34352
rect 10875 34318 10909 34352
rect 10943 34318 10977 34352
rect 11011 34318 11045 34352
rect 11079 34318 11113 34352
rect 11147 34318 11181 34352
rect 11215 34318 11249 34352
rect 11283 34318 11317 34352
rect 11351 34318 11385 34352
rect 11419 34318 11453 34352
rect 11487 34318 11521 34352
rect 11555 34318 11589 34352
rect 11623 34318 11657 34352
rect 11691 34328 11781 34352
rect 11854 34350 11912 34424
rect 12850 34350 12920 34424
rect 12992 34351 13062 34424
rect 16100 34352 16192 34424
rect 15203 34351 15227 34352
rect 11691 34318 11747 34328
rect 9445 34278 9479 34318
rect 9445 34210 9479 34244
rect 11747 34260 11781 34294
rect 11747 34192 11781 34226
rect 11374 34187 11747 34188
rect 9445 34142 9479 34176
rect 9445 34098 9479 34108
rect 9775 34181 10321 34187
rect 9775 34147 9836 34181
rect 9870 34147 9970 34181
rect 10004 34147 10092 34181
rect 10126 34147 10226 34181
rect 10260 34147 10321 34181
rect 9775 34141 10321 34147
rect 9657 34098 9711 34099
rect 9445 34074 9711 34098
rect 9479 34068 9711 34074
rect 9479 34040 9667 34068
rect 9445 34020 9667 34040
rect 9701 34020 9711 34068
rect 9445 34006 9711 34020
rect 9479 33996 9711 34006
rect 9479 33972 9667 33996
rect 9445 33938 9479 33972
rect 9445 33870 9479 33904
rect 9445 33802 9479 33836
rect 9445 33734 9479 33768
rect 9445 33666 9479 33700
rect 8583 33644 8659 33663
rect 7892 33610 7926 33644
rect 6986 33585 7342 33592
rect 6952 33551 7342 33585
rect 6986 33536 7342 33551
rect 6952 33483 6986 33517
rect 7142 33473 7342 33536
rect 7892 33542 7926 33576
rect 7892 33474 7926 33508
rect 6952 33415 6986 33449
rect 7604 33387 7650 33414
rect 7892 33406 7926 33440
rect 6952 33347 6986 33381
rect 7342 33353 7650 33387
rect 7692 33353 7802 33387
rect 6952 33279 6986 33313
rect 7892 33338 7926 33372
rect 8034 33634 8438 33644
rect 8034 33600 8317 33634
rect 8351 33600 8438 33634
rect 8034 33584 8438 33600
rect 8583 33610 8606 33644
rect 8640 33610 8659 33644
rect 8583 33591 8659 33610
rect 9445 33598 9479 33632
rect 8034 33388 8094 33584
rect 8245 33493 8300 33547
rect 8248 33406 8282 33493
rect 8456 33400 8490 33546
rect 8664 33418 8698 33496
rect 8729 33493 8784 33547
rect 8944 33436 8978 33543
rect 8940 33402 8978 33436
rect 9445 33530 9479 33564
rect 9657 33952 9667 33972
rect 9701 33952 9711 33996
rect 9657 33924 9711 33952
rect 9657 33884 9667 33924
rect 9701 33884 9711 33924
rect 9657 33852 9711 33884
rect 9657 33816 9667 33852
rect 9701 33816 9711 33852
rect 9657 33782 9711 33816
rect 9657 33746 9667 33782
rect 9701 33746 9711 33782
rect 9657 33714 9711 33746
rect 9657 33674 9667 33714
rect 9701 33674 9711 33714
rect 9657 33646 9711 33674
rect 9657 33602 9667 33646
rect 9701 33602 9711 33646
rect 9657 33578 9711 33602
rect 9657 33530 9667 33578
rect 9701 33530 9711 33578
rect 9657 33499 9711 33530
rect 9775 34054 9809 34141
rect 9775 33986 9809 34020
rect 9775 33918 9809 33952
rect 9775 33850 9809 33884
rect 9775 33782 9809 33816
rect 9775 33714 9809 33748
rect 9775 33646 9809 33680
rect 9775 33578 9809 33612
rect 9445 33462 9479 33496
rect 8034 33354 8045 33388
rect 8079 33354 8094 33388
rect 8034 33340 8094 33354
rect 9445 33394 9479 33428
rect 9775 33457 9809 33544
rect 10031 34054 10065 34141
rect 10031 33986 10065 34020
rect 10031 33918 10065 33952
rect 10031 33850 10065 33884
rect 10031 33782 10065 33816
rect 10031 33714 10065 33748
rect 10031 33646 10065 33680
rect 10031 33578 10065 33612
rect 10031 33457 10065 33544
rect 10287 34054 10321 34141
rect 10905 34181 11747 34187
rect 10905 34147 10966 34181
rect 11000 34147 11100 34181
rect 11134 34147 11222 34181
rect 11256 34147 11356 34181
rect 11390 34158 11747 34181
rect 11390 34147 11781 34158
rect 10905 34141 11781 34147
rect 10287 33986 10321 34020
rect 10287 33918 10321 33952
rect 10287 33850 10321 33884
rect 10287 33782 10321 33816
rect 10287 33714 10321 33748
rect 10287 33646 10321 33680
rect 10287 33578 10321 33612
rect 10287 33499 10321 33544
rect 10543 34054 10577 34099
rect 10543 33986 10577 34020
rect 10543 33918 10577 33952
rect 10543 33850 10577 33884
rect 10543 33782 10577 33816
rect 10543 33714 10577 33748
rect 10543 33646 10577 33680
rect 10543 33578 10577 33612
rect 10543 33457 10577 33544
rect 10649 34054 10683 34099
rect 10649 33986 10683 34020
rect 10649 33918 10683 33952
rect 10649 33850 10683 33884
rect 10649 33782 10683 33816
rect 10649 33714 10683 33748
rect 10649 33646 10683 33680
rect 10649 33578 10683 33612
rect 10649 33499 10683 33544
rect 10905 34054 10939 34141
rect 10905 33986 10939 34020
rect 10905 33918 10939 33952
rect 10905 33850 10939 33884
rect 10905 33782 10939 33816
rect 10905 33714 10939 33748
rect 10905 33646 10939 33680
rect 10905 33578 10939 33612
rect 10905 33499 10939 33544
rect 11161 34054 11195 34141
rect 11374 34140 11781 34141
rect 11161 33986 11195 34020
rect 11161 33918 11195 33952
rect 11161 33850 11195 33884
rect 11161 33782 11195 33816
rect 11161 33714 11195 33748
rect 11161 33646 11195 33680
rect 11161 33578 11195 33612
rect 11161 33499 11195 33544
rect 11417 34054 11451 34140
rect 11747 34124 11781 34140
rect 11417 33986 11451 34020
rect 11417 33918 11451 33952
rect 11417 33850 11451 33884
rect 11417 33782 11451 33816
rect 11417 33714 11451 33748
rect 11417 33646 11451 33680
rect 11417 33578 11451 33612
rect 11417 33457 11451 33544
rect 11515 34068 11569 34099
rect 11515 34020 11525 34068
rect 11559 34020 11569 34068
rect 11515 33996 11569 34020
rect 11515 33952 11525 33996
rect 11559 33952 11569 33996
rect 11515 33924 11569 33952
rect 11515 33884 11525 33924
rect 11559 33884 11569 33924
rect 11515 33852 11569 33884
rect 11515 33816 11525 33852
rect 11559 33816 11569 33852
rect 11515 33782 11569 33816
rect 11515 33746 11525 33782
rect 11559 33746 11569 33782
rect 11515 33714 11569 33746
rect 11515 33674 11525 33714
rect 11559 33674 11569 33714
rect 11515 33646 11569 33674
rect 11515 33602 11525 33646
rect 11559 33602 11569 33646
rect 11515 33578 11569 33602
rect 11515 33530 11525 33578
rect 11559 33530 11569 33578
rect 11515 33499 11569 33530
rect 11747 34056 11781 34090
rect 11747 33988 11781 34022
rect 11747 33920 11781 33954
rect 11747 33852 11781 33886
rect 11747 33784 11781 33818
rect 11747 33716 11781 33750
rect 11747 33648 11781 33682
rect 11747 33580 11781 33614
rect 11747 33512 11781 33546
rect 9775 33451 10276 33457
rect 9775 33417 9836 33451
rect 9870 33417 9970 33451
rect 10004 33417 10092 33451
rect 10126 33417 10226 33451
rect 10260 33417 10276 33451
rect 9775 33411 10276 33417
rect 10332 33451 10577 33457
rect 10332 33417 10348 33451
rect 10382 33417 10482 33451
rect 10516 33417 10577 33451
rect 10332 33411 10577 33417
rect 10694 33451 10894 33457
rect 10694 33417 10710 33451
rect 10744 33417 10844 33451
rect 10878 33417 10894 33451
rect 10694 33411 10894 33417
rect 10950 33451 11150 33457
rect 10950 33417 10966 33451
rect 11000 33417 11100 33451
rect 11134 33417 11150 33451
rect 10950 33411 11150 33417
rect 11206 33451 11451 33457
rect 11206 33417 11222 33451
rect 11256 33417 11356 33451
rect 11390 33417 11451 33451
rect 11206 33411 11451 33417
rect 11747 33444 11781 33478
rect 7892 33255 7926 33304
rect 9445 33326 9479 33360
rect 9445 33258 9479 33292
rect 6986 33245 7052 33255
rect 6952 33221 7052 33245
rect 7086 33221 7120 33255
rect 7154 33221 7188 33255
rect 7222 33221 7256 33255
rect 7290 33221 7324 33255
rect 7358 33221 7392 33255
rect 7426 33221 7460 33255
rect 7494 33221 7528 33255
rect 7562 33221 7596 33255
rect 7630 33221 7664 33255
rect 7698 33221 7732 33255
rect 7766 33221 7800 33255
rect 7834 33221 7868 33255
rect 7902 33221 7926 33255
rect 7514 33176 7562 33178
rect 8074 33176 8122 33194
rect 7514 33172 8122 33176
rect 7514 33138 7521 33172
rect 7555 33171 8122 33172
rect 7555 33138 8078 33171
rect 7514 33137 8078 33138
rect 8112 33137 8122 33171
rect 8162 33183 8196 33223
rect 8334 33186 8368 33223
rect 8334 33183 8506 33186
rect 8162 33172 8506 33183
rect 8162 33149 8446 33172
rect 7514 33132 8122 33137
rect 7514 33130 7562 33132
rect 8074 33116 8122 33132
rect 8334 33138 8446 33149
rect 8480 33138 8506 33172
rect 8334 33126 8506 33138
rect 7638 33092 7662 33098
rect 6952 33058 6976 33092
rect 7010 33058 7044 33092
rect 7078 33058 7112 33092
rect 7146 33058 7180 33092
rect 7214 33058 7248 33092
rect 7282 33058 7316 33092
rect 7350 33058 7384 33092
rect 7418 33058 7452 33092
rect 7486 33058 7520 33092
rect 7554 33064 7662 33092
rect 7696 33064 7730 33098
rect 7764 33064 7798 33098
rect 7832 33092 7924 33098
rect 7832 33064 7914 33092
rect 7554 33058 7672 33064
rect 7890 33058 7914 33064
rect 7948 33058 8036 33092
rect 8334 33091 8368 33126
rect 6952 32976 6986 33058
rect 8002 33040 8036 33058
rect 8320 33057 8368 33091
rect 8542 33057 8576 33238
rect 8822 33186 8856 33241
rect 8822 33174 8988 33186
rect 8736 33170 8988 33174
rect 8736 33136 8926 33170
rect 8960 33136 8988 33170
rect 8736 33126 8988 33136
rect 9029 33184 9063 33257
rect 11747 33376 11781 33410
rect 11747 33308 11781 33342
rect 11747 33234 11781 33274
rect 9479 33224 9547 33234
rect 9445 33200 9547 33224
rect 9581 33200 9615 33234
rect 9649 33200 9683 33234
rect 9717 33200 9751 33234
rect 9785 33200 9819 33234
rect 9853 33200 9887 33234
rect 9921 33200 9955 33234
rect 9989 33200 10023 33234
rect 10057 33200 10091 33234
rect 10125 33200 10159 33234
rect 10193 33200 10227 33234
rect 10261 33200 10295 33234
rect 10329 33200 10363 33234
rect 10397 33200 10431 33234
rect 10465 33200 10499 33234
rect 10533 33200 10567 33234
rect 10601 33200 10635 33234
rect 10669 33200 10703 33234
rect 10737 33200 10771 33234
rect 10805 33200 10839 33234
rect 10873 33200 10907 33234
rect 10941 33200 10975 33234
rect 11009 33200 11043 33234
rect 11077 33200 11111 33234
rect 11145 33200 11179 33234
rect 11213 33200 11247 33234
rect 11281 33200 11315 33234
rect 11349 33200 11383 33234
rect 11417 33200 11451 33234
rect 11485 33200 11519 33234
rect 11553 33200 11587 33234
rect 11621 33200 11655 33234
rect 11689 33200 11723 33234
rect 11757 33200 11781 33234
rect 11853 34316 11877 34350
rect 11911 34316 11945 34350
rect 11979 34316 12013 34350
rect 12047 34316 12081 34350
rect 12115 34316 12149 34350
rect 12183 34316 12217 34350
rect 12251 34316 12285 34350
rect 12319 34316 12353 34350
rect 12387 34316 12421 34350
rect 12455 34316 12489 34350
rect 12523 34316 12557 34350
rect 12591 34316 12625 34350
rect 12659 34316 12693 34350
rect 12727 34316 12761 34350
rect 12795 34334 12920 34350
rect 12795 34326 12919 34334
rect 12795 34316 12885 34326
rect 11853 34248 11887 34316
rect 12885 34258 12919 34292
rect 11853 34241 12885 34248
rect 11887 34238 12885 34241
rect 11887 34207 11998 34238
rect 11853 34204 11998 34207
rect 12036 34204 12070 34238
rect 12104 34204 12138 34238
rect 12176 34204 12258 34238
rect 12296 34204 12330 34238
rect 12364 34204 12398 34238
rect 12436 34204 12499 34238
rect 12539 34204 12571 34238
rect 12607 34204 12641 34238
rect 12677 34204 12709 34238
rect 12749 34224 12885 34238
rect 12991 34317 13015 34351
rect 13049 34317 13083 34351
rect 13117 34317 13151 34351
rect 13185 34317 13219 34351
rect 13253 34317 13287 34351
rect 13321 34317 13355 34351
rect 13389 34317 13423 34351
rect 13457 34317 13491 34351
rect 13525 34317 13559 34351
rect 13593 34317 13627 34351
rect 13661 34317 13695 34351
rect 13729 34317 13763 34351
rect 13797 34317 13831 34351
rect 13865 34317 13899 34351
rect 13933 34317 13967 34351
rect 14001 34317 14035 34351
rect 14069 34317 14103 34351
rect 14137 34317 14171 34351
rect 14205 34317 14239 34351
rect 14273 34317 14307 34351
rect 14341 34317 14375 34351
rect 14409 34317 14443 34351
rect 14477 34317 14511 34351
rect 14545 34317 14579 34351
rect 14613 34317 14647 34351
rect 14681 34317 14715 34351
rect 14749 34317 14783 34351
rect 14817 34317 14851 34351
rect 14885 34317 14919 34351
rect 14953 34317 14987 34351
rect 15021 34317 15055 34351
rect 15089 34317 15123 34351
rect 15157 34318 15227 34351
rect 15261 34318 15295 34352
rect 15329 34318 15363 34352
rect 15397 34318 15431 34352
rect 15465 34318 15499 34352
rect 15533 34318 15567 34352
rect 15601 34318 15635 34352
rect 15669 34318 15703 34352
rect 15737 34318 15771 34352
rect 15805 34318 15839 34352
rect 15873 34318 15907 34352
rect 15941 34318 15975 34352
rect 16009 34318 16043 34352
rect 16077 34328 16193 34352
rect 16077 34318 16159 34328
rect 15157 34317 15237 34318
rect 12991 34278 13025 34317
rect 12919 34244 12991 34248
rect 16159 34260 16193 34294
rect 13025 34244 13026 34248
rect 12919 34230 13026 34244
rect 12919 34224 15781 34230
rect 12749 34220 15781 34224
rect 12749 34210 13119 34220
rect 12749 34204 12991 34210
rect 11853 34194 12991 34204
rect 11853 34173 11887 34194
rect 11853 34105 11887 34139
rect 11853 34037 11887 34071
rect 11853 33969 11887 34003
rect 11853 33901 11887 33935
rect 11853 33833 11887 33867
rect 11853 33734 11887 33799
rect 11853 33666 11887 33700
rect 11853 33598 11887 33632
rect 11853 33530 11887 33564
rect 11853 33462 11887 33496
rect 11853 33394 11887 33428
rect 11963 34092 11997 34194
rect 11963 34024 11997 34058
rect 11963 33956 11997 33990
rect 11963 33888 11997 33922
rect 11963 33820 11997 33854
rect 11963 33752 11997 33786
rect 11963 33684 11997 33718
rect 11963 33616 11997 33650
rect 11963 33548 11997 33582
rect 11963 33480 11997 33514
rect 11963 33414 11997 33446
rect 12219 34092 12253 34124
rect 12219 34024 12253 34058
rect 12219 33956 12253 33990
rect 12219 33888 12253 33922
rect 12219 33820 12253 33854
rect 12219 33752 12253 33786
rect 12219 33684 12253 33718
rect 12219 33616 12253 33650
rect 12219 33548 12253 33582
rect 12219 33480 12253 33514
rect 12219 33414 12253 33446
rect 12475 34092 12509 34194
rect 12874 34190 12991 34194
rect 12874 34176 12885 34190
rect 12919 34176 12991 34190
rect 13025 34186 13119 34210
rect 13171 34186 13187 34220
rect 13243 34186 13255 34220
rect 13315 34186 13323 34220
rect 13387 34186 13391 34220
rect 13493 34186 13497 34220
rect 13561 34186 13569 34220
rect 13629 34186 13641 34220
rect 13697 34186 13713 34220
rect 13765 34186 13893 34220
rect 13945 34186 13961 34220
rect 14017 34186 14029 34220
rect 14089 34186 14097 34220
rect 14161 34186 14165 34220
rect 14267 34186 14271 34220
rect 14335 34186 14343 34220
rect 14403 34186 14415 34220
rect 14471 34186 14487 34220
rect 14539 34186 15781 34220
rect 13025 34176 15781 34186
rect 15880 34226 16159 34230
rect 15880 34192 16193 34226
rect 15880 34176 16159 34192
rect 12475 34024 12509 34058
rect 12475 33956 12509 33990
rect 12475 33888 12509 33922
rect 12475 33820 12509 33854
rect 12475 33752 12509 33786
rect 12475 33684 12509 33718
rect 12475 33616 12509 33650
rect 12475 33548 12509 33582
rect 12475 33480 12509 33514
rect 12475 33414 12509 33446
rect 12731 34092 12765 34124
rect 12731 34024 12765 34058
rect 12731 33956 12765 33990
rect 12731 33888 12765 33922
rect 12731 33820 12765 33854
rect 12731 33752 12765 33786
rect 12731 33684 12765 33718
rect 12731 33616 12765 33650
rect 12731 33548 12765 33582
rect 12731 33480 12765 33514
rect 12731 33414 12765 33446
rect 12885 34122 12919 34156
rect 12885 34054 12919 34088
rect 12885 33986 12919 34020
rect 12885 33918 12919 33952
rect 12885 33850 12919 33884
rect 12885 33782 12919 33816
rect 12885 33714 12919 33748
rect 12885 33646 12919 33680
rect 12885 33578 12919 33612
rect 12885 33510 12919 33544
rect 12885 33442 12919 33476
rect 12885 33374 12919 33408
rect 11853 33326 11887 33360
rect 12008 33366 12208 33372
rect 12008 33332 12024 33366
rect 12058 33332 12158 33366
rect 12192 33332 12208 33366
rect 12008 33326 12208 33332
rect 12264 33366 12464 33372
rect 12264 33332 12280 33366
rect 12314 33332 12414 33366
rect 12448 33332 12464 33366
rect 12264 33326 12464 33332
rect 12520 33366 12720 33372
rect 12520 33332 12536 33366
rect 12570 33332 12670 33366
rect 12704 33332 12720 33366
rect 12520 33326 12720 33332
rect 11853 33258 11887 33292
rect 12885 33306 12919 33340
rect 12885 33234 12919 33272
rect 11887 33224 11977 33234
rect 11853 33200 11977 33224
rect 12011 33200 12045 33234
rect 12079 33200 12113 33234
rect 12147 33200 12181 33234
rect 12215 33200 12249 33234
rect 12283 33200 12317 33234
rect 12351 33200 12385 33234
rect 12419 33200 12453 33234
rect 12487 33200 12521 33234
rect 12555 33200 12589 33234
rect 12623 33200 12657 33234
rect 12691 33200 12725 33234
rect 12759 33200 12793 33234
rect 12827 33200 12861 33234
rect 12895 33200 12919 33234
rect 12991 34142 13025 34176
rect 12991 34074 13025 34108
rect 12991 34006 13025 34040
rect 12991 33938 13025 33972
rect 12991 33870 13025 33904
rect 12991 33802 13025 33836
rect 12991 33734 13025 33768
rect 12991 33666 13025 33700
rect 12991 33598 13025 33632
rect 12991 33530 13025 33564
rect 12991 33462 13025 33496
rect 12991 33394 13025 33428
rect 12991 33326 13025 33360
rect 13097 34057 13131 34176
rect 13097 33989 13131 34023
rect 13097 33921 13131 33955
rect 13097 33853 13131 33887
rect 13097 33785 13131 33819
rect 13097 33717 13131 33751
rect 13097 33649 13131 33683
rect 13097 33581 13131 33615
rect 13097 33513 13131 33547
rect 13097 33389 13131 33479
rect 13753 34057 13787 34176
rect 13753 33989 13787 34023
rect 13753 33921 13787 33955
rect 13753 33853 13787 33887
rect 13753 33785 13787 33819
rect 13753 33717 13787 33751
rect 13753 33649 13787 33683
rect 13753 33581 13787 33615
rect 13753 33513 13787 33547
rect 13753 33389 13787 33479
rect 13875 34057 13909 34106
rect 13875 33989 13909 34023
rect 13875 33921 13909 33955
rect 13875 33853 13909 33887
rect 13875 33785 13909 33819
rect 13875 33717 13909 33751
rect 13875 33649 13909 33683
rect 13875 33581 13909 33615
rect 13875 33513 13909 33547
rect 13875 33431 13909 33479
rect 14531 34057 14565 34176
rect 15309 34106 15343 34176
rect 15965 34106 15999 34176
rect 16159 34124 16193 34158
rect 14531 33989 14565 34023
rect 14531 33921 14565 33955
rect 14531 33853 14565 33887
rect 14531 33785 14565 33819
rect 14531 33717 14565 33751
rect 14531 33649 14565 33683
rect 14531 33581 14565 33615
rect 14531 33513 14565 33547
rect 14531 33431 14565 33479
rect 16159 34056 16193 34090
rect 16159 33988 16193 34022
rect 19229 33993 19340 34193
rect 19392 33993 19426 34193
rect 16159 33920 16193 33954
rect 16159 33852 16193 33886
rect 19330 33882 19400 33902
rect 19330 33848 19348 33882
rect 19382 33848 19400 33882
rect 19330 33830 19400 33848
rect 16159 33784 16193 33818
rect 16159 33716 16193 33750
rect 16159 33648 16193 33682
rect 16159 33580 16193 33614
rect 16159 33512 16193 33546
rect 16159 33444 16193 33478
rect 15187 33389 15221 33431
rect 13097 33383 13787 33389
rect 13097 33349 13158 33383
rect 13192 33349 13234 33383
rect 13268 33349 13310 33383
rect 13344 33349 13386 33383
rect 13420 33349 13462 33383
rect 13496 33349 13538 33383
rect 13572 33349 13615 33383
rect 13649 33349 13692 33383
rect 13726 33349 13787 33383
rect 13097 33343 13787 33349
rect 13920 33383 14520 33389
rect 13920 33349 13936 33383
rect 13970 33349 14012 33383
rect 14046 33349 14088 33383
rect 14122 33349 14164 33383
rect 14198 33349 14240 33383
rect 14274 33349 14316 33383
rect 14350 33349 14393 33383
rect 14427 33349 14470 33383
rect 14504 33349 14520 33383
rect 13920 33343 14520 33349
rect 15157 33343 15221 33389
rect 15309 33389 15343 33431
rect 15965 33389 15999 33431
rect 15309 33343 15429 33389
rect 15919 33343 15999 33389
rect 16159 33376 16193 33410
rect 12991 33258 13025 33292
rect 16159 33308 16193 33342
rect 16159 33234 16193 33274
rect 13025 33224 13106 33234
rect 12991 33200 13106 33224
rect 13140 33200 13174 33234
rect 13208 33200 13242 33234
rect 13276 33200 13310 33234
rect 13344 33200 13378 33234
rect 13412 33200 13446 33234
rect 13480 33200 13514 33234
rect 13548 33200 13582 33234
rect 13616 33200 13650 33234
rect 13684 33200 13718 33234
rect 13752 33200 13786 33234
rect 13820 33200 13854 33234
rect 13888 33200 13922 33234
rect 13956 33200 13990 33234
rect 14024 33200 14058 33234
rect 14092 33200 14126 33234
rect 14160 33200 14194 33234
rect 14228 33200 14262 33234
rect 14296 33200 14330 33234
rect 14364 33200 14398 33234
rect 14432 33200 14466 33234
rect 14500 33200 14534 33234
rect 14568 33200 14639 33234
rect 14673 33200 14707 33234
rect 14741 33200 14775 33234
rect 14809 33200 14843 33234
rect 14877 33200 14911 33234
rect 14945 33200 14979 33234
rect 15013 33200 15047 33234
rect 15081 33200 15115 33234
rect 15149 33200 15183 33234
rect 15217 33200 15251 33234
rect 15285 33200 15319 33234
rect 15353 33200 15387 33234
rect 15421 33200 15455 33234
rect 15489 33200 15523 33234
rect 15557 33200 15591 33234
rect 15625 33200 15659 33234
rect 15693 33200 15727 33234
rect 15761 33200 15795 33234
rect 15829 33200 15863 33234
rect 15897 33200 15931 33234
rect 15965 33200 15999 33234
rect 16033 33200 16067 33234
rect 16101 33200 16135 33234
rect 16169 33200 16193 33234
rect 9029 33170 9146 33184
rect 9029 33136 9096 33170
rect 9130 33136 9146 33170
rect 8736 33091 8770 33126
rect 9029 33120 9146 33136
rect 9029 33058 9063 33120
rect 7366 32993 7446 33024
rect 8002 33016 8072 33040
rect 8002 33006 8038 33016
rect 6952 32908 6986 32942
rect 7142 32934 7242 32968
rect 7366 32959 7389 32993
rect 7423 32959 7446 32993
rect 7366 32934 7446 32959
rect 7570 32970 7948 33004
rect 7570 32903 7604 32970
rect 7742 32908 7776 32970
rect 7914 32915 7948 32970
rect 8038 32948 8072 32982
rect 9434 33004 9458 33038
rect 9492 33004 9526 33038
rect 9560 33004 9594 33038
rect 9628 33004 9662 33038
rect 9696 33004 9730 33038
rect 9764 33004 9798 33038
rect 9832 33004 9866 33038
rect 9900 33004 9934 33038
rect 9968 33004 10002 33038
rect 10036 33004 10070 33038
rect 10104 33004 10138 33038
rect 10172 33004 10206 33038
rect 10240 33004 10274 33038
rect 10308 33004 10342 33038
rect 10376 33004 10410 33038
rect 10444 33004 10478 33038
rect 10512 33004 10546 33038
rect 10580 33004 10614 33038
rect 10648 33004 10682 33038
rect 10716 33004 10750 33038
rect 10784 33004 10818 33038
rect 10852 33004 10886 33038
rect 10920 33004 10954 33038
rect 10988 33004 11022 33038
rect 11056 33004 11090 33038
rect 11124 33004 11158 33038
rect 11192 33014 11422 33038
rect 11192 33004 11242 33014
rect 6952 32840 6986 32874
rect 6952 32772 6986 32806
rect 6952 32704 6986 32738
rect 6952 32636 6986 32670
rect 6952 32568 6986 32602
rect 6952 32500 6986 32534
rect 6952 32432 6986 32466
rect 6952 32364 6986 32398
rect 6952 32296 6986 32330
rect 6952 32228 6986 32262
rect 6952 32160 6986 32194
rect 6952 32092 6986 32126
rect 6952 32024 6986 32058
rect 6952 31956 6986 31990
rect 6854 31898 6878 31932
rect 6912 31922 6952 31932
rect 6912 31898 6986 31922
rect 8038 32880 8072 32914
rect 8530 32946 8590 32960
rect 8530 32912 8542 32946
rect 8576 32912 8590 32946
rect 9434 32927 9468 33004
rect 8038 32822 8072 32846
rect 8162 32822 8196 32891
rect 8456 32822 8490 32898
rect 8530 32894 8590 32912
rect 8650 32822 8684 32906
rect 8822 32822 8856 32913
rect 8943 32822 8977 32915
rect 11276 33004 11330 33014
rect 11242 32946 11276 32980
rect 9468 32910 11093 32920
rect 9468 32893 9642 32910
rect 9434 32876 9642 32893
rect 9684 32876 9714 32910
rect 9752 32876 9786 32910
rect 9820 32876 9854 32910
rect 9892 32876 9922 32910
rect 9964 32876 10038 32910
rect 10078 32876 10110 32910
rect 10146 32876 10180 32910
rect 10216 32876 10248 32910
rect 10288 32876 10394 32910
rect 10434 32876 10466 32910
rect 10502 32876 10536 32910
rect 10572 32876 10604 32910
rect 10644 32876 10735 32910
rect 10777 32876 10807 32910
rect 10845 32876 10879 32910
rect 10913 32876 10947 32910
rect 10985 32876 11015 32910
rect 11057 32876 11093 32910
rect 9434 32866 11093 32876
rect 11364 33004 11422 33014
rect 11456 33004 11490 33038
rect 11524 33004 11558 33038
rect 11592 33004 11626 33038
rect 11660 33004 11694 33038
rect 11728 33004 11762 33038
rect 11796 33004 11830 33038
rect 11864 33004 11898 33038
rect 11932 33004 11966 33038
rect 12000 33004 12034 33038
rect 12068 33004 12102 33038
rect 12136 33004 12170 33038
rect 12204 33004 12238 33038
rect 12272 33004 12306 33038
rect 12340 33004 12374 33038
rect 12408 33004 12442 33038
rect 12476 33004 12510 33038
rect 12544 33004 12578 33038
rect 12612 33004 12646 33038
rect 12680 33004 12714 33038
rect 12748 33004 12782 33038
rect 12816 33004 12850 33038
rect 12884 33004 12918 33038
rect 12952 33004 12986 33038
rect 13020 33004 13054 33038
rect 13088 33004 13122 33038
rect 13156 33004 13190 33038
rect 13224 33004 13258 33038
rect 13292 33004 13326 33038
rect 13360 33004 13394 33038
rect 13428 33004 13462 33038
rect 13496 33004 13530 33038
rect 13564 33004 13598 33038
rect 13632 33004 13666 33038
rect 13700 33004 13734 33038
rect 13768 33004 13802 33038
rect 13836 33004 13870 33038
rect 13904 33004 13938 33038
rect 13972 33004 14006 33038
rect 14040 33004 14074 33038
rect 14108 33004 14142 33038
rect 14176 33004 14210 33038
rect 14244 33004 14278 33038
rect 14312 33004 14346 33038
rect 14380 33004 14414 33038
rect 14448 33004 14482 33038
rect 14516 33004 14550 33038
rect 14584 33004 14618 33038
rect 14652 33004 14686 33038
rect 14720 33004 14754 33038
rect 14788 33004 14822 33038
rect 14856 33004 14890 33038
rect 14924 33004 14958 33038
rect 14992 33004 15026 33038
rect 15060 33004 15094 33038
rect 15128 33004 15162 33038
rect 15196 33004 15230 33038
rect 15264 33004 15298 33038
rect 15332 33004 15366 33038
rect 15400 33004 15434 33038
rect 15468 33004 15502 33038
rect 15536 33004 15570 33038
rect 15604 33004 15638 33038
rect 15672 33004 15706 33038
rect 15740 33004 15774 33038
rect 15808 33004 15842 33038
rect 15876 33004 15910 33038
rect 15944 33004 15978 33038
rect 16012 33004 16046 33038
rect 16080 33004 16114 33038
rect 16148 33004 16182 33038
rect 16216 33004 16250 33038
rect 16284 33004 16318 33038
rect 16352 33004 16376 33038
rect 11330 32946 11364 32980
rect 11242 32878 11276 32912
rect 11326 32912 11330 32936
rect 16342 32970 16376 33004
rect 11364 32930 11995 32936
rect 11364 32912 11511 32930
rect 11326 32896 11511 32912
rect 11545 32896 11584 32930
rect 11618 32896 11657 32930
rect 11691 32896 11729 32930
rect 11763 32896 11801 32930
rect 11835 32896 11873 32930
rect 11907 32896 11945 32930
rect 11979 32896 11995 32930
rect 11326 32890 11995 32896
rect 12051 32930 12551 32936
rect 12051 32896 12067 32930
rect 12101 32896 12140 32930
rect 12174 32896 12213 32930
rect 12247 32896 12285 32930
rect 12319 32896 12357 32930
rect 12391 32896 12429 32930
rect 12463 32896 12501 32930
rect 12535 32896 12551 32930
rect 12051 32890 12551 32896
rect 12607 32930 13107 32936
rect 12607 32896 12623 32930
rect 12657 32896 12695 32930
rect 12729 32896 12767 32930
rect 12801 32896 12839 32930
rect 12873 32896 12911 32930
rect 12945 32896 12984 32930
rect 13018 32896 13057 32930
rect 13091 32896 13107 32930
rect 12607 32890 13107 32896
rect 13224 32930 13769 32936
rect 13224 32896 13285 32930
rect 13319 32896 13357 32930
rect 13391 32896 13429 32930
rect 13463 32896 13501 32930
rect 13535 32896 13573 32930
rect 13607 32896 13646 32930
rect 13680 32896 13719 32930
rect 13753 32896 13769 32930
rect 13224 32890 13769 32896
rect 13825 32930 14391 32936
rect 13825 32896 13841 32930
rect 13875 32896 13914 32930
rect 13948 32896 13987 32930
rect 14021 32896 14059 32930
rect 14093 32896 14131 32930
rect 14165 32896 14203 32930
rect 14237 32896 14275 32930
rect 14309 32896 14391 32930
rect 13825 32890 14391 32896
rect 16186 32902 16376 32936
rect 16186 32890 16342 32902
rect 9434 32859 9468 32866
rect 9434 32822 9468 32825
rect 8038 32812 9468 32822
rect 8072 32791 9468 32812
rect 11242 32810 11276 32844
rect 8072 32778 9434 32791
rect 8038 32762 9434 32778
rect 8038 32744 8072 32762
rect 8038 32676 8072 32710
rect 8870 32710 8938 32726
rect 8870 32676 8886 32710
rect 8920 32676 8938 32710
rect 8870 32656 8938 32676
rect 9434 32723 9468 32757
rect 8038 32608 8072 32642
rect 8038 32540 8072 32574
rect 8038 32472 8072 32506
rect 8038 32404 8072 32438
rect 8038 32336 8072 32370
rect 8038 32268 8072 32302
rect 8038 32200 8072 32234
rect 8038 32132 8072 32166
rect 8038 32064 8072 32098
rect 8038 31963 8072 32030
rect 6854 31827 6888 31898
rect 8038 31895 8072 31929
rect 6854 31759 6888 31793
rect 6854 31691 6888 31725
rect 6854 31623 6888 31657
rect 7142 31599 7242 31888
rect 8038 31827 8072 31861
rect 8038 31759 8072 31793
rect 8038 31691 8072 31725
rect 8038 31623 8072 31657
rect 6888 31589 6928 31599
rect 6854 31565 6928 31589
rect 6962 31565 6996 31599
rect 7030 31565 7064 31599
rect 7098 31565 7132 31599
rect 7166 31565 7200 31599
rect 7234 31565 7268 31599
rect 7302 31565 7336 31599
rect 7370 31565 7394 31599
rect 7360 31468 7394 31565
rect 7360 31400 7394 31434
rect 7360 31332 7394 31366
rect 7360 31264 7394 31298
rect 7360 31196 7394 31230
rect 7360 31128 7394 31162
rect 7360 31060 7394 31094
rect 7360 30992 7394 31026
rect 7331 30958 7360 30968
rect 8038 31555 8072 31589
rect 8038 31487 8072 31521
rect 8038 31419 8072 31453
rect 8038 31351 8072 31385
rect 8038 31283 8072 31317
rect 8038 31215 8072 31249
rect 8038 31147 8072 31181
rect 8038 31079 8072 31113
rect 8038 30968 8072 31045
rect 9434 32655 9468 32689
rect 9434 32587 9468 32621
rect 9434 32519 9468 32553
rect 9434 32451 9468 32485
rect 9434 32383 9468 32417
rect 9434 32315 9468 32349
rect 9434 32247 9468 32281
rect 9434 32179 9468 32213
rect 9434 32111 9468 32145
rect 9434 32043 9468 32077
rect 9434 31975 9468 32009
rect 9434 31907 9468 31941
rect 9434 31839 9468 31873
rect 9434 31771 9468 31805
rect 9434 31703 9468 31737
rect 9434 31635 9468 31669
rect 9434 31567 9468 31601
rect 9434 31499 9468 31533
rect 9434 31431 9468 31465
rect 9434 31363 9468 31397
rect 9629 32757 9663 32794
rect 9629 32689 9663 32723
rect 9629 32621 9663 32655
rect 9629 32553 9663 32587
rect 9629 32485 9663 32519
rect 9629 32417 9663 32451
rect 9629 32349 9663 32383
rect 9629 32281 9663 32315
rect 9629 32213 9663 32247
rect 9629 32145 9663 32179
rect 9629 32077 9663 32111
rect 9629 32009 9663 32043
rect 9629 31941 9663 31975
rect 9629 31873 9663 31907
rect 9629 31805 9663 31839
rect 9629 31737 9663 31771
rect 9629 31669 9663 31703
rect 9629 31601 9663 31635
rect 9629 31533 9663 31567
rect 9629 31465 9663 31499
rect 9629 31394 9663 31431
rect 9985 32757 10019 32794
rect 9985 32689 10019 32723
rect 9985 32621 10019 32655
rect 9985 32553 10019 32587
rect 9985 32485 10019 32519
rect 9985 32417 10019 32451
rect 9985 32349 10019 32383
rect 9985 32281 10019 32315
rect 9985 32213 10019 32247
rect 9985 32145 10019 32179
rect 9985 32077 10019 32111
rect 9985 32009 10019 32043
rect 9985 31941 10019 31975
rect 9985 31873 10019 31907
rect 9985 31805 10019 31839
rect 9985 31737 10019 31771
rect 9985 31669 10019 31703
rect 9985 31601 10019 31635
rect 9985 31533 10019 31567
rect 9985 31465 10019 31499
rect 9985 31394 10019 31431
rect 10341 32757 10375 32794
rect 10341 32689 10375 32723
rect 10341 32621 10375 32655
rect 10341 32553 10375 32587
rect 10341 32485 10375 32519
rect 10341 32417 10375 32451
rect 10341 32349 10375 32383
rect 10341 32281 10375 32315
rect 10341 32213 10375 32247
rect 10341 32145 10375 32179
rect 10341 32077 10375 32111
rect 10341 32009 10375 32043
rect 10341 31941 10375 31975
rect 10341 31873 10375 31907
rect 10341 31805 10375 31839
rect 10341 31737 10375 31771
rect 10341 31669 10375 31703
rect 10341 31601 10375 31635
rect 10341 31533 10375 31567
rect 10341 31465 10375 31499
rect 10341 31394 10375 31431
rect 10697 32757 10731 32794
rect 10697 32689 10731 32723
rect 10697 32621 10731 32655
rect 10697 32553 10731 32587
rect 10697 32485 10731 32519
rect 10697 32417 10731 32451
rect 10697 32349 10731 32383
rect 10697 32281 10731 32315
rect 10697 32213 10731 32247
rect 10697 32145 10731 32179
rect 10697 32077 10731 32111
rect 10697 32009 10731 32043
rect 10697 31941 10731 31975
rect 10697 31873 10731 31907
rect 10697 31805 10731 31839
rect 10697 31737 10731 31771
rect 10697 31669 10731 31703
rect 10697 31601 10731 31635
rect 10697 31533 10731 31567
rect 10697 31465 10731 31499
rect 10697 31394 10731 31431
rect 11053 32757 11087 32794
rect 11053 32689 11087 32723
rect 11053 32621 11087 32655
rect 11242 32742 11276 32776
rect 11242 32674 11276 32708
rect 11242 32606 11276 32640
rect 11087 32587 11138 32590
rect 11053 32578 11138 32587
rect 11053 32553 11091 32578
rect 11087 32544 11091 32553
rect 11125 32544 11138 32578
rect 11087 32530 11138 32544
rect 11242 32538 11276 32572
rect 11053 32485 11087 32519
rect 11053 32417 11087 32451
rect 11053 32349 11087 32383
rect 11053 32281 11087 32315
rect 11053 32213 11087 32247
rect 11053 32145 11087 32179
rect 11053 32077 11087 32111
rect 11053 32009 11087 32043
rect 11053 31941 11087 31975
rect 11053 31873 11087 31907
rect 11053 31805 11087 31839
rect 11053 31737 11087 31771
rect 11053 31669 11087 31703
rect 11053 31601 11087 31635
rect 11053 31533 11087 31567
rect 11053 31465 11087 31499
rect 11053 31394 11087 31431
rect 11242 32470 11276 32504
rect 11242 32402 11276 32436
rect 11242 32334 11276 32368
rect 11242 32266 11276 32300
rect 11242 32198 11276 32232
rect 11242 32130 11276 32164
rect 11242 32062 11276 32096
rect 11242 31994 11276 32028
rect 11242 31926 11276 31960
rect 11242 31858 11276 31892
rect 11242 31790 11276 31824
rect 11242 31722 11276 31756
rect 11242 31654 11276 31688
rect 11242 31586 11276 31620
rect 11330 32878 11364 32890
rect 11330 32810 11364 32844
rect 11330 32742 11364 32776
rect 11330 32674 11364 32708
rect 11330 32606 11364 32640
rect 11330 32538 11364 32572
rect 11330 32470 11364 32504
rect 11330 32402 11364 32436
rect 11330 32334 11364 32368
rect 11330 32266 11364 32300
rect 11330 32198 11364 32232
rect 11330 32130 11364 32164
rect 11330 32062 11364 32096
rect 11330 31994 11364 32028
rect 11330 31926 11364 31960
rect 11330 31858 11364 31892
rect 11330 31790 11364 31824
rect 11330 31722 11364 31756
rect 11450 32819 11484 32890
rect 11450 32751 11484 32785
rect 11450 32683 11484 32717
rect 11450 32615 11484 32649
rect 11450 32547 11484 32581
rect 11450 32479 11484 32513
rect 11450 32411 11484 32445
rect 11450 32265 11484 32377
rect 11450 32197 11484 32231
rect 11450 32129 11484 32163
rect 11450 32061 11484 32095
rect 11450 31993 11484 32027
rect 11450 31925 11484 31959
rect 11450 31857 11484 31891
rect 11450 31722 11484 31823
rect 12006 32819 12040 32848
rect 12006 32751 12040 32785
rect 12006 32683 12040 32717
rect 12006 32615 12040 32649
rect 12006 32547 12040 32581
rect 12006 32479 12040 32513
rect 12006 32411 12040 32445
rect 12006 32265 12040 32377
rect 12006 32197 12040 32231
rect 12006 32129 12040 32163
rect 12006 32061 12040 32095
rect 12006 31993 12040 32027
rect 12006 31925 12040 31959
rect 12006 31857 12040 31891
rect 12006 31722 12040 31823
rect 12562 32819 12596 32848
rect 12562 32751 12596 32785
rect 12562 32683 12596 32717
rect 12562 32615 12596 32649
rect 12562 32547 12596 32581
rect 12562 32479 12596 32513
rect 12562 32411 12596 32445
rect 12562 32265 12596 32377
rect 12562 32197 12596 32231
rect 12562 32129 12596 32163
rect 12562 32061 12596 32095
rect 12562 31993 12596 32027
rect 12562 31925 12596 31959
rect 12562 31857 12596 31891
rect 12562 31794 12596 31823
rect 13118 32819 13152 32848
rect 13118 32751 13152 32785
rect 13118 32683 13152 32717
rect 13118 32615 13152 32649
rect 13118 32547 13152 32581
rect 13118 32479 13152 32513
rect 13118 32411 13152 32445
rect 13118 32265 13152 32377
rect 13118 32197 13152 32231
rect 13118 32129 13152 32163
rect 13118 32061 13152 32095
rect 13118 31993 13152 32027
rect 13118 31925 13152 31959
rect 13118 31857 13152 31891
rect 13118 31722 13152 31823
rect 13224 32819 13258 32890
rect 13224 32751 13258 32785
rect 13224 32683 13258 32717
rect 13224 32615 13258 32649
rect 13224 32547 13258 32581
rect 13224 32479 13258 32513
rect 13224 32411 13258 32445
rect 13224 32265 13258 32377
rect 13224 32197 13258 32231
rect 13224 32129 13258 32163
rect 13224 32061 13258 32095
rect 13224 31993 13258 32027
rect 13224 31925 13258 31959
rect 13224 31857 13258 31891
rect 13224 31794 13258 31823
rect 13780 32819 13814 32848
rect 13780 32751 13814 32785
rect 13780 32683 13814 32717
rect 13780 32615 13814 32649
rect 13780 32547 13814 32581
rect 13780 32479 13814 32513
rect 13780 32411 13814 32445
rect 13780 32265 13814 32377
rect 13780 32197 13814 32231
rect 13780 32129 13814 32163
rect 13780 32061 13814 32095
rect 13780 31993 13814 32027
rect 13780 31925 13814 31959
rect 13780 31857 13814 31891
rect 13780 31722 13814 31823
rect 14336 32819 14370 32890
rect 16214 32848 16248 32890
rect 14336 32751 14370 32785
rect 14336 32683 14370 32717
rect 14336 32615 14370 32649
rect 14336 32547 14370 32581
rect 14336 32479 14370 32513
rect 14336 32411 14370 32445
rect 16342 32834 16376 32868
rect 16342 32766 16376 32800
rect 16342 32698 16376 32732
rect 16342 32630 16376 32664
rect 16342 32562 16376 32596
rect 16342 32494 16376 32528
rect 16342 32426 16376 32460
rect 14336 32265 14370 32377
rect 14440 32268 14474 32348
rect 14996 32252 15030 32348
rect 15102 32263 15136 32382
rect 16342 32358 16376 32392
rect 15658 32262 15692 32352
rect 16214 32262 16248 32352
rect 16342 32290 16376 32324
rect 14336 32197 14370 32231
rect 14336 32129 14370 32163
rect 14336 32061 14370 32095
rect 14336 31993 14370 32027
rect 14336 31925 14370 31959
rect 14336 31857 14370 31891
rect 14336 31794 14370 31823
rect 16342 32222 16376 32256
rect 16342 32154 16376 32188
rect 16342 32086 16376 32120
rect 16342 32018 16376 32052
rect 16342 31950 16376 31984
rect 16342 31882 16376 31916
rect 16342 31814 16376 31848
rect 14440 31722 14474 31796
rect 15658 31722 15692 31796
rect 16214 31722 16248 31796
rect 16342 31746 16376 31780
rect 11364 31712 14485 31722
rect 11364 31688 11469 31712
rect 11330 31678 11469 31688
rect 11525 31678 11537 31712
rect 11597 31678 11605 31712
rect 11669 31678 11673 31712
rect 11775 31678 11779 31712
rect 11843 31678 11851 31712
rect 11911 31678 11923 31712
rect 11979 31678 12051 31712
rect 12097 31678 12123 31712
rect 12165 31678 12195 31712
rect 12233 31678 12267 31712
rect 12301 31678 12335 31712
rect 12373 31678 12403 31712
rect 12445 31678 12471 31712
rect 12517 31678 12592 31712
rect 12640 31678 12664 31712
rect 12708 31678 12736 31712
rect 12776 31678 12808 31712
rect 12844 31678 12878 31712
rect 12914 31678 12946 31712
rect 12986 31678 13014 31712
rect 13058 31678 13082 31712
rect 13130 31678 13246 31712
rect 13294 31678 13318 31712
rect 13362 31678 13390 31712
rect 13430 31678 13462 31712
rect 13498 31678 13532 31712
rect 13568 31678 13600 31712
rect 13640 31678 13668 31712
rect 13712 31678 13736 31712
rect 13784 31678 13841 31712
rect 13897 31678 13909 31712
rect 13969 31678 13977 31712
rect 14041 31678 14045 31712
rect 14147 31678 14151 31712
rect 14215 31678 14223 31712
rect 14283 31678 14295 31712
rect 14351 31678 14485 31712
rect 11330 31668 14485 31678
rect 14992 31668 15154 31722
rect 15607 31668 15769 31722
rect 16198 31712 16342 31722
rect 16198 31678 16376 31712
rect 16198 31668 16342 31678
rect 11330 31654 11364 31668
rect 11330 31586 11364 31620
rect 16342 31610 16376 31644
rect 12668 31586 14656 31588
rect 11276 31552 11354 31586
rect 11388 31552 11422 31586
rect 11456 31552 11490 31586
rect 11524 31552 11558 31586
rect 11592 31552 11626 31586
rect 11660 31552 11694 31586
rect 11728 31552 11762 31586
rect 11796 31552 11830 31586
rect 11864 31552 11898 31586
rect 11932 31552 11966 31586
rect 12000 31552 12034 31586
rect 12068 31552 12102 31586
rect 12136 31552 12170 31586
rect 12204 31552 12238 31586
rect 12272 31552 12306 31586
rect 12340 31552 12374 31586
rect 12408 31552 12442 31586
rect 12476 31552 12510 31586
rect 12544 31552 12578 31586
rect 12612 31552 12646 31586
rect 12680 31552 12714 31586
rect 12748 31552 12782 31586
rect 12816 31552 12850 31586
rect 12884 31552 12918 31586
rect 12952 31552 12986 31586
rect 13020 31552 13054 31586
rect 13088 31552 13122 31586
rect 13156 31552 13190 31586
rect 13224 31552 13258 31586
rect 13292 31552 13326 31586
rect 13360 31552 13394 31586
rect 13428 31552 13462 31586
rect 13496 31552 13530 31586
rect 13564 31552 13598 31586
rect 13632 31552 13666 31586
rect 13700 31552 13734 31586
rect 13768 31552 13877 31586
rect 13911 31552 13945 31586
rect 13979 31552 14013 31586
rect 14047 31552 14081 31586
rect 14115 31552 14149 31586
rect 14183 31552 14217 31586
rect 14251 31552 14285 31586
rect 14319 31552 14353 31586
rect 14387 31552 14421 31586
rect 14455 31552 14489 31586
rect 14523 31552 14557 31586
rect 14591 31552 14625 31586
rect 14659 31552 14693 31586
rect 14727 31552 14761 31586
rect 14795 31552 14829 31586
rect 14863 31552 14897 31586
rect 14931 31552 14965 31586
rect 14999 31552 15033 31586
rect 15067 31552 15101 31586
rect 15135 31552 15169 31586
rect 15203 31552 15237 31586
rect 15271 31552 15305 31586
rect 15339 31552 15373 31586
rect 15407 31552 15441 31586
rect 15475 31552 15509 31586
rect 15543 31552 15577 31586
rect 15611 31552 15645 31586
rect 15679 31552 15713 31586
rect 15747 31552 15781 31586
rect 15815 31552 15849 31586
rect 15883 31552 15917 31586
rect 15951 31552 15985 31586
rect 16019 31552 16053 31586
rect 16087 31552 16121 31586
rect 16155 31552 16189 31586
rect 16223 31552 16257 31586
rect 16291 31576 16342 31586
rect 16291 31552 16376 31576
rect 11242 31518 11276 31552
rect 11242 31450 11276 31484
rect 11242 31382 11276 31416
rect 9434 31295 9468 31329
rect 9674 31346 9974 31352
rect 9674 31312 9690 31346
rect 9724 31312 9768 31346
rect 9802 31312 9846 31346
rect 9880 31312 9924 31346
rect 9958 31312 9974 31346
rect 9674 31306 9974 31312
rect 10030 31346 10330 31352
rect 10030 31312 10046 31346
rect 10080 31312 10124 31346
rect 10158 31312 10202 31346
rect 10236 31312 10280 31346
rect 10314 31312 10330 31346
rect 10030 31306 10330 31312
rect 10386 31346 10686 31352
rect 10386 31312 10402 31346
rect 10436 31312 10480 31346
rect 10514 31312 10558 31346
rect 10592 31312 10636 31346
rect 10670 31312 10686 31346
rect 10386 31306 10686 31312
rect 10742 31346 11042 31352
rect 10742 31312 10758 31346
rect 10792 31312 10836 31346
rect 10870 31312 10914 31346
rect 10948 31312 10992 31346
rect 11026 31312 11042 31346
rect 10742 31306 11042 31312
rect 11522 31351 11722 31552
rect 12668 31380 14656 31552
rect 11242 31314 11276 31348
rect 9434 31194 9468 31261
rect 11242 31246 11276 31280
rect 12668 31346 12777 31380
rect 12811 31346 12845 31380
rect 12879 31346 12913 31380
rect 12947 31346 12981 31380
rect 13015 31346 13049 31380
rect 13083 31346 13117 31380
rect 13151 31346 13185 31380
rect 13219 31346 13253 31380
rect 13287 31346 13321 31380
rect 13355 31346 13389 31380
rect 13423 31346 13457 31380
rect 13491 31346 13525 31380
rect 13559 31346 13593 31380
rect 13627 31346 13661 31380
rect 13695 31346 13729 31380
rect 13763 31346 13797 31380
rect 13831 31346 13865 31380
rect 13899 31346 13933 31380
rect 13967 31346 14001 31380
rect 14035 31346 14069 31380
rect 14103 31346 14137 31380
rect 14171 31346 14205 31380
rect 14239 31346 14273 31380
rect 14307 31346 14341 31380
rect 14375 31346 14409 31380
rect 14443 31346 14477 31380
rect 14511 31348 14656 31380
rect 14511 31346 14620 31348
rect 12668 31266 12702 31346
rect 11242 31178 11276 31212
rect 9434 31126 9468 31160
rect 9674 31162 9974 31168
rect 9674 31128 9690 31162
rect 9724 31128 9768 31162
rect 9802 31128 9846 31162
rect 9880 31128 9924 31162
rect 9958 31128 9974 31162
rect 9674 31122 9974 31128
rect 10030 31162 10330 31168
rect 10030 31128 10046 31162
rect 10080 31128 10124 31162
rect 10158 31128 10202 31162
rect 10236 31128 10280 31162
rect 10314 31128 10330 31162
rect 10030 31122 10330 31128
rect 10386 31162 10686 31168
rect 10386 31128 10402 31162
rect 10436 31128 10480 31162
rect 10514 31128 10558 31162
rect 10592 31128 10636 31162
rect 10670 31128 10686 31162
rect 10386 31122 10686 31128
rect 10742 31162 11042 31168
rect 10742 31128 10758 31162
rect 10792 31128 10836 31162
rect 10870 31128 10914 31162
rect 10948 31128 10992 31162
rect 11026 31128 11042 31162
rect 10742 31122 11042 31128
rect 9434 31058 9468 31092
rect 11242 31110 11276 31144
rect 11376 31190 11446 31206
rect 11655 31199 11883 31233
rect 14586 31266 14620 31346
rect 11376 31156 11396 31190
rect 11430 31156 11446 31190
rect 11376 31138 11446 31156
rect 12668 31198 12702 31232
rect 14586 31198 14620 31232
rect 9434 30990 9468 31024
rect 7331 30934 7394 30958
rect 7331 30850 7365 30934
rect 7484 30850 7518 30930
rect 7656 30850 7690 30961
rect 8038 30944 8101 30968
rect 8038 30934 8067 30944
rect 7828 30850 7862 30922
rect 8067 30876 8101 30910
rect 7331 30843 8067 30850
rect 7365 30842 8067 30843
rect 7365 30809 8101 30842
rect 7331 30808 8101 30809
rect 7331 30796 8067 30808
rect 7331 30775 7365 30796
rect 7331 30707 7365 30741
rect 8067 30683 8101 30774
rect 7365 30673 7431 30683
rect 7331 30649 7431 30673
rect 7465 30649 7499 30683
rect 7533 30649 7567 30683
rect 7601 30649 7635 30683
rect 7669 30649 7703 30683
rect 7737 30649 7771 30683
rect 7805 30649 7839 30683
rect 7873 30649 7907 30683
rect 7941 30649 7975 30683
rect 8009 30649 8043 30683
rect 8077 30649 8101 30683
rect 9434 30922 9468 30956
rect 9434 30854 9468 30888
rect 9434 30786 9468 30820
rect 9434 30718 9468 30752
rect 9434 30650 9468 30684
rect 9434 30582 9468 30616
rect 9434 30514 9468 30548
rect 9434 30446 9468 30480
rect 9434 30378 9468 30412
rect 9434 30310 9468 30344
rect 9434 30242 9468 30276
rect 9434 30174 9468 30208
rect 9434 30106 9468 30140
rect 9434 30038 9468 30072
rect 9434 29970 9468 30004
rect 9434 29902 9468 29936
rect 9434 29834 9468 29868
rect 9434 29766 9468 29800
rect 9434 29698 9468 29732
rect 9629 31043 9663 31080
rect 9629 30975 9663 31009
rect 9629 30907 9663 30941
rect 9629 30839 9663 30873
rect 9629 30771 9663 30805
rect 9629 30703 9663 30737
rect 9629 30635 9663 30669
rect 9629 30567 9663 30601
rect 9629 30499 9663 30533
rect 9629 30431 9663 30465
rect 9629 30363 9663 30397
rect 9629 30295 9663 30329
rect 9629 30227 9663 30261
rect 9629 30159 9663 30193
rect 9985 31043 10019 31080
rect 9985 30975 10019 31009
rect 9985 30907 10019 30941
rect 9985 30839 10019 30873
rect 9985 30771 10019 30805
rect 9985 30703 10019 30737
rect 9985 30635 10019 30669
rect 9985 30567 10019 30601
rect 9985 30499 10019 30533
rect 9985 30431 10019 30465
rect 9985 30363 10019 30397
rect 9985 30295 10019 30329
rect 9985 30227 10019 30261
rect 9985 30159 10019 30193
rect 9629 30091 9663 30125
rect 9629 30023 9663 30057
rect 9629 29955 9663 29989
rect 9629 29887 9663 29921
rect 9629 29819 9663 29853
rect 9984 30104 9985 30154
rect 10341 31043 10375 31080
rect 10341 30975 10375 31009
rect 10341 30907 10375 30941
rect 10341 30839 10375 30873
rect 10341 30771 10375 30805
rect 10341 30703 10375 30737
rect 10341 30635 10375 30669
rect 10341 30567 10375 30601
rect 10341 30499 10375 30533
rect 10341 30431 10375 30465
rect 10341 30363 10375 30397
rect 10341 30295 10375 30329
rect 10341 30227 10375 30261
rect 10341 30159 10375 30193
rect 10019 30104 10020 30154
rect 9984 30091 10020 30104
rect 9984 30032 9985 30091
rect 10019 30032 10020 30091
rect 9984 30023 10020 30032
rect 9984 29960 9985 30023
rect 10019 29960 10020 30023
rect 9984 29955 10020 29960
rect 9984 29888 9985 29955
rect 10019 29888 10020 29955
rect 9984 29887 10020 29888
rect 9984 29853 9985 29887
rect 10019 29853 10020 29887
rect 9984 29850 10020 29853
rect 9984 29800 9985 29850
rect 9629 29751 9663 29785
rect 9629 29680 9663 29717
rect 10019 29800 10020 29850
rect 10341 30091 10375 30125
rect 10341 30023 10375 30057
rect 10341 29955 10375 29989
rect 10341 29887 10375 29921
rect 10341 29819 10375 29853
rect 9985 29751 10019 29785
rect 9985 29680 10019 29717
rect 10341 29751 10375 29785
rect 10341 29680 10375 29717
rect 10697 31043 10731 31080
rect 10697 30975 10731 31009
rect 10697 30907 10731 30941
rect 10697 30839 10731 30873
rect 10697 30771 10731 30805
rect 10697 30703 10731 30737
rect 10697 30635 10731 30669
rect 10697 30567 10731 30601
rect 10697 30499 10731 30533
rect 10697 30431 10731 30465
rect 10697 30363 10731 30397
rect 10697 30295 10731 30329
rect 10697 30227 10731 30261
rect 10697 30159 10731 30193
rect 10697 30091 10731 30125
rect 10697 30023 10731 30057
rect 10697 29955 10731 29989
rect 10697 29887 10731 29921
rect 10697 29819 10731 29853
rect 10697 29751 10731 29785
rect 10697 29680 10731 29717
rect 11053 31043 11087 31080
rect 11053 30975 11087 31009
rect 11053 30907 11087 30941
rect 11053 30839 11087 30873
rect 11053 30771 11087 30805
rect 11053 30703 11087 30737
rect 11053 30635 11087 30669
rect 11053 30567 11087 30601
rect 11053 30499 11087 30533
rect 11053 30431 11087 30465
rect 11053 30363 11087 30397
rect 11053 30295 11087 30329
rect 11053 30227 11087 30261
rect 11053 30159 11087 30193
rect 11053 30091 11087 30125
rect 11053 30023 11087 30057
rect 11053 29955 11087 29989
rect 11053 29887 11087 29921
rect 11053 29819 11087 29853
rect 11053 29751 11087 29785
rect 11053 29680 11087 29717
rect 11242 31042 11276 31076
rect 12668 31084 12702 31164
rect 14586 31084 14620 31164
rect 12668 31050 12777 31084
rect 12811 31050 12845 31084
rect 12879 31050 12913 31084
rect 12947 31050 12981 31084
rect 13015 31050 13049 31084
rect 13083 31050 13117 31084
rect 13151 31050 13185 31084
rect 13219 31050 13253 31084
rect 13287 31050 13321 31084
rect 13355 31050 13389 31084
rect 13423 31050 13457 31084
rect 13491 31050 13525 31084
rect 13559 31050 13593 31084
rect 13627 31050 13661 31084
rect 13695 31050 13729 31084
rect 13763 31050 13797 31084
rect 13831 31050 13865 31084
rect 13899 31050 13933 31084
rect 13967 31050 14001 31084
rect 14035 31050 14069 31084
rect 14103 31050 14137 31084
rect 14171 31050 14205 31084
rect 14239 31050 14273 31084
rect 14307 31050 14341 31084
rect 14375 31050 14409 31084
rect 14443 31050 14477 31084
rect 14511 31050 14620 31084
rect 11242 30974 11276 31008
rect 11242 30906 11276 30940
rect 11242 30838 11276 30872
rect 11242 30770 11276 30804
rect 11242 30702 11276 30736
rect 11242 30634 11276 30668
rect 11242 30566 11276 30600
rect 11242 30498 11276 30532
rect 11242 30430 11276 30464
rect 11242 30362 11276 30396
rect 11242 30294 11276 30328
rect 11242 30226 11276 30260
rect 11242 30158 11276 30192
rect 11242 30090 11276 30124
rect 11242 30022 11276 30056
rect 11242 29954 11276 29988
rect 11242 29886 11276 29920
rect 11242 29818 11276 29852
rect 11242 29750 11276 29784
rect 11242 29682 11276 29716
rect 9434 29630 9468 29664
rect 11242 29614 11276 29648
rect 9468 29598 11242 29608
rect 9468 29596 9659 29598
rect 9434 29564 9659 29596
rect 9701 29564 9731 29598
rect 9769 29564 9803 29598
rect 9837 29564 9871 29598
rect 9909 29564 9939 29598
rect 9981 29564 10072 29598
rect 10112 29564 10144 29598
rect 10180 29564 10214 29598
rect 10250 29564 10282 29598
rect 10322 29564 10411 29598
rect 10451 29564 10483 29598
rect 10519 29564 10553 29598
rect 10589 29564 10621 29598
rect 10661 29564 10735 29598
rect 10777 29564 10807 29598
rect 10845 29564 10879 29598
rect 10913 29564 10947 29598
rect 10985 29564 11015 29598
rect 11057 29580 11242 29598
rect 11057 29564 11276 29580
rect 9434 29562 11276 29564
rect 9468 29554 11276 29562
rect 9434 29494 9468 29528
rect 11242 29546 11276 29554
rect 11242 29470 11276 29512
rect 9468 29460 9518 29470
rect 9434 29436 9518 29460
rect 9552 29436 9586 29470
rect 9620 29436 9654 29470
rect 9688 29436 9722 29470
rect 9756 29436 9790 29470
rect 9824 29436 9858 29470
rect 9892 29436 9926 29470
rect 9960 29436 9994 29470
rect 10028 29436 10062 29470
rect 10096 29436 10130 29470
rect 10164 29436 10198 29470
rect 10232 29436 10266 29470
rect 10300 29436 10334 29470
rect 10368 29436 10402 29470
rect 10436 29436 10470 29470
rect 10504 29436 10538 29470
rect 10572 29436 10606 29470
rect 10640 29436 10674 29470
rect 10708 29436 10742 29470
rect 10776 29436 10810 29470
rect 10844 29436 10878 29470
rect 10912 29436 10946 29470
rect 10980 29436 11014 29470
rect 11048 29436 11082 29470
rect 11116 29436 11150 29470
rect 11184 29436 11218 29470
rect 11252 29436 11276 29470
rect 9434 28480 9640 29436
rect 12236 28874 12858 29306
rect 8236 25776 8306 27516
rect 8634 25766 8704 27588
rect 9524 25760 9594 27582
rect 9922 25766 9992 27588
rect 10814 25766 10884 27588
rect 12236 27434 12518 28448
rect 12236 26576 12858 27008
rect 10962 25148 11768 25580
rect 13326 24812 13608 25580
rect 10924 24712 13608 24812
rect 11457 19226 11481 19260
rect 11515 19226 11549 19260
rect 11583 19226 11617 19260
rect 11651 19226 11685 19260
rect 11719 19226 11753 19260
rect 11787 19226 11821 19260
rect 11855 19226 11889 19260
rect 11923 19226 11957 19260
rect 11991 19226 12025 19260
rect 12059 19226 12093 19260
rect 12127 19226 12161 19260
rect 12195 19226 12229 19260
rect 12263 19226 12297 19260
rect 12331 19226 12365 19260
rect 12399 19226 12433 19260
rect 12467 19226 12501 19260
rect 12535 19226 12569 19260
rect 12603 19226 12637 19260
rect 12671 19226 12705 19260
rect 12739 19226 12773 19260
rect 12807 19226 12841 19260
rect 12875 19226 12909 19260
rect 12943 19226 12977 19260
rect 13011 19226 13045 19260
rect 13079 19226 13113 19260
rect 13147 19226 13181 19260
rect 13215 19226 13249 19260
rect 13283 19226 13317 19260
rect 13351 19226 13385 19260
rect 13419 19226 13453 19260
rect 13487 19226 13521 19260
rect 13555 19226 13589 19260
rect 13623 19226 13657 19260
rect 13691 19226 13725 19260
rect 13759 19226 13793 19260
rect 13827 19226 13861 19260
rect 13895 19226 13929 19260
rect 13963 19226 13997 19260
rect 14031 19226 14065 19260
rect 14099 19226 14133 19260
rect 14167 19226 14201 19260
rect 14235 19226 14269 19260
rect 14303 19226 14360 19260
rect 14394 19226 14428 19260
rect 14462 19226 14496 19260
rect 14530 19226 14564 19260
rect 14598 19226 14632 19260
rect 14666 19226 14700 19260
rect 14734 19226 14768 19260
rect 14802 19226 14836 19260
rect 14870 19226 14904 19260
rect 14938 19226 14972 19260
rect 15006 19226 15040 19260
rect 15074 19226 15108 19260
rect 15142 19226 15176 19260
rect 15210 19226 15244 19260
rect 15278 19226 15312 19260
rect 15346 19226 15380 19260
rect 15414 19226 15448 19260
rect 15482 19226 15516 19260
rect 15550 19226 15584 19260
rect 15618 19226 15652 19260
rect 15686 19226 15720 19260
rect 15754 19226 15788 19260
rect 15822 19226 15856 19260
rect 15890 19226 15924 19260
rect 15958 19226 15992 19260
rect 16026 19226 16060 19260
rect 16094 19226 16128 19260
rect 16162 19226 16196 19260
rect 16230 19226 16264 19260
rect 16298 19226 16332 19260
rect 16366 19226 16400 19260
rect 16434 19226 16468 19260
rect 16502 19226 16536 19260
rect 16570 19226 16604 19260
rect 16638 19226 16672 19260
rect 16706 19226 16740 19260
rect 16774 19226 16808 19260
rect 16842 19226 16876 19260
rect 16910 19226 16944 19260
rect 16978 19226 17012 19260
rect 17046 19226 17080 19260
rect 17114 19236 17383 19260
rect 17114 19226 17181 19236
rect 11457 19166 11491 19226
rect 17215 19202 17287 19236
rect 17321 19226 17383 19236
rect 17417 19226 17451 19260
rect 17485 19226 17519 19260
rect 17553 19226 17587 19260
rect 17621 19226 17655 19260
rect 17689 19226 17723 19260
rect 17757 19226 17791 19260
rect 17825 19226 17859 19260
rect 17893 19226 17927 19260
rect 17961 19226 17995 19260
rect 18029 19226 18063 19260
rect 18097 19226 18131 19260
rect 18165 19226 18199 19260
rect 18233 19226 18267 19260
rect 18301 19226 18335 19260
rect 18369 19226 18403 19260
rect 18437 19226 18471 19260
rect 18505 19226 18539 19260
rect 18573 19226 18607 19260
rect 18641 19226 18675 19260
rect 18709 19226 18743 19260
rect 18777 19226 18811 19260
rect 18845 19226 18879 19260
rect 18913 19226 18947 19260
rect 18981 19226 19015 19260
rect 19049 19226 19083 19260
rect 19117 19226 19151 19260
rect 19185 19226 19219 19260
rect 19253 19226 19287 19260
rect 19321 19226 19355 19260
rect 19389 19226 19423 19260
rect 19457 19226 19491 19260
rect 19525 19226 19559 19260
rect 19593 19226 19627 19260
rect 19661 19226 19695 19260
rect 19729 19226 19763 19260
rect 19797 19226 19831 19260
rect 19865 19226 19899 19260
rect 19933 19226 19967 19260
rect 20001 19226 20035 19260
rect 20069 19226 20103 19260
rect 20137 19226 20171 19260
rect 20205 19236 20374 19260
rect 20205 19226 20301 19236
rect 17181 19168 17321 19202
rect 17215 19134 17287 19168
rect 11491 19132 11583 19134
rect 11457 19098 11583 19132
rect 11491 19080 11583 19098
rect 12279 19080 12389 19134
rect 12953 19080 13063 19134
rect 13590 19080 13700 19134
rect 14264 19080 14374 19134
rect 14950 19080 15060 19134
rect 15610 19080 15720 19134
rect 16303 19080 16413 19134
rect 17084 19116 17321 19134
rect 20195 19202 20301 19226
rect 20335 19226 20374 19236
rect 20408 19226 20442 19260
rect 20476 19226 20510 19260
rect 20544 19226 20578 19260
rect 20612 19226 20646 19260
rect 20680 19226 20714 19260
rect 20748 19226 20782 19260
rect 20816 19226 20850 19260
rect 20884 19226 20918 19260
rect 20952 19226 20986 19260
rect 21020 19226 21054 19260
rect 21088 19226 21122 19260
rect 21156 19226 21190 19260
rect 21224 19226 21258 19260
rect 21292 19226 21326 19260
rect 21360 19226 21394 19260
rect 21428 19226 21462 19260
rect 21496 19226 21530 19260
rect 21564 19226 21598 19260
rect 21632 19226 21666 19260
rect 21700 19226 21734 19260
rect 21768 19226 21802 19260
rect 21836 19226 21870 19260
rect 21904 19226 21938 19260
rect 21972 19226 22006 19260
rect 22040 19226 22074 19260
rect 22108 19226 22142 19260
rect 22176 19226 22210 19260
rect 22244 19226 22278 19260
rect 22312 19226 22346 19260
rect 22380 19226 22414 19260
rect 22448 19226 22482 19260
rect 22516 19226 22550 19260
rect 22584 19226 22618 19260
rect 22652 19226 22686 19260
rect 22720 19226 22754 19260
rect 22788 19226 22822 19260
rect 22856 19226 22890 19260
rect 22924 19226 22958 19260
rect 22992 19226 23026 19260
rect 23060 19226 23157 19260
rect 23191 19226 23225 19260
rect 23259 19226 23293 19260
rect 23327 19226 23361 19260
rect 23395 19226 23429 19260
rect 23463 19226 23497 19260
rect 23531 19226 23565 19260
rect 23599 19226 23633 19260
rect 23667 19226 23701 19260
rect 23735 19226 23769 19260
rect 23803 19226 23837 19260
rect 23871 19226 23905 19260
rect 23939 19226 23973 19260
rect 24007 19226 24041 19260
rect 24075 19226 24109 19260
rect 24143 19226 24177 19260
rect 24211 19226 24245 19260
rect 24279 19226 24313 19260
rect 24347 19226 24381 19260
rect 24415 19226 24449 19260
rect 24483 19226 24517 19260
rect 24551 19226 24585 19260
rect 24619 19226 24653 19260
rect 24687 19226 24721 19260
rect 24755 19226 24789 19260
rect 24823 19226 24857 19260
rect 24891 19226 24925 19260
rect 24959 19226 24993 19260
rect 25027 19226 25061 19260
rect 25095 19226 25129 19260
rect 25163 19226 25197 19260
rect 25231 19226 25265 19260
rect 25299 19226 25333 19260
rect 25367 19226 25401 19260
rect 25435 19226 25469 19260
rect 25503 19226 25537 19260
rect 25571 19226 25605 19260
rect 25639 19226 25673 19260
rect 25707 19226 25741 19260
rect 25775 19226 25809 19260
rect 25843 19226 25867 19260
rect 20195 19168 20335 19202
rect 20195 19140 20301 19168
rect 17084 19100 17428 19116
rect 17084 19080 17181 19100
rect 11457 19030 11491 19064
rect 13662 19006 13698 19080
rect 14974 19004 15010 19080
rect 17215 19066 17287 19100
rect 17321 19066 17428 19100
rect 17181 19062 17428 19066
rect 18035 19062 18145 19116
rect 18703 19062 18813 19116
rect 19397 19062 19507 19116
rect 20089 19106 20195 19116
rect 20229 19134 20301 19140
rect 20229 19116 20335 19134
rect 25833 19166 25867 19226
rect 25833 19116 25867 19132
rect 20229 19106 20444 19116
rect 20089 19100 20444 19106
rect 20089 19072 20301 19100
rect 20089 19062 20195 19072
rect 17181 19032 17321 19062
rect 11457 18962 11491 18996
rect 11457 18894 11491 18928
rect 11457 18826 11491 18860
rect 11457 18758 11491 18792
rect 11457 18690 11491 18724
rect 11457 18622 11491 18656
rect 11457 18554 11491 18588
rect 11457 18486 11491 18520
rect 11457 18418 11491 18452
rect 11457 18350 11491 18384
rect 11457 18282 11491 18316
rect 11457 18214 11491 18248
rect 11457 18146 11491 18180
rect 11457 18078 11491 18112
rect 11457 18010 11491 18044
rect 11457 17942 11491 17976
rect 11457 17874 11491 17908
rect 11457 17806 11491 17840
rect 11457 17738 11491 17772
rect 11457 17670 11491 17704
rect 17215 18998 17287 19032
rect 17181 18964 17321 18998
rect 18740 18988 18776 19062
rect 20229 19066 20301 19072
rect 20335 19066 20444 19100
rect 20229 19062 20444 19066
rect 21054 19062 21164 19116
rect 21735 19062 21845 19116
rect 22368 19062 22478 19116
rect 23035 19062 23145 19116
rect 23669 19062 23779 19116
rect 24353 19062 24463 19116
rect 25033 19062 25143 19116
rect 25727 19098 25867 19116
rect 25727 19064 25833 19098
rect 25727 19062 25867 19064
rect 20229 19038 20335 19062
rect 20195 19032 20335 19038
rect 20195 19004 20301 19032
rect 17215 18930 17287 18964
rect 17181 18896 17321 18930
rect 17215 18862 17287 18896
rect 17181 18828 17321 18862
rect 17215 18794 17287 18828
rect 17181 18760 17321 18794
rect 17215 18726 17287 18760
rect 17181 18692 17321 18726
rect 17215 18658 17287 18692
rect 17181 18624 17321 18658
rect 17215 18590 17287 18624
rect 17181 18556 17321 18590
rect 17215 18522 17287 18556
rect 17181 18488 17321 18522
rect 17215 18454 17287 18488
rect 17181 18420 17321 18454
rect 17215 18386 17287 18420
rect 17181 18352 17321 18386
rect 17215 18318 17287 18352
rect 17181 18284 17321 18318
rect 17215 18250 17287 18284
rect 17181 18216 17321 18250
rect 17215 18182 17287 18216
rect 17181 18148 17321 18182
rect 17215 18114 17287 18148
rect 17181 18080 17321 18114
rect 17215 18046 17287 18080
rect 17181 18012 17321 18046
rect 17215 17978 17287 18012
rect 17181 17944 17321 17978
rect 17215 17910 17287 17944
rect 17181 17876 17321 17910
rect 17215 17842 17287 17876
rect 17181 17808 17321 17842
rect 17215 17774 17287 17808
rect 17181 17740 17321 17774
rect 17215 17706 17287 17740
rect 20229 18998 20301 19004
rect 20229 18970 20335 18998
rect 21755 18979 21789 19062
rect 23722 18982 23758 19062
rect 25034 18978 25070 19062
rect 25833 19030 25867 19062
rect 20195 18964 20335 18970
rect 20195 18936 20301 18964
rect 20229 18930 20301 18936
rect 20229 18902 20335 18930
rect 20195 18896 20335 18902
rect 20195 18868 20301 18896
rect 20229 18862 20301 18868
rect 20229 18834 20335 18862
rect 20195 18828 20335 18834
rect 20195 18800 20301 18828
rect 20229 18794 20301 18800
rect 20229 18766 20335 18794
rect 20195 18760 20335 18766
rect 20195 18732 20301 18760
rect 20229 18726 20301 18732
rect 20229 18698 20335 18726
rect 20195 18692 20335 18698
rect 20195 18664 20301 18692
rect 20229 18658 20301 18664
rect 20229 18630 20335 18658
rect 20195 18624 20335 18630
rect 20195 18596 20301 18624
rect 20229 18590 20301 18596
rect 20229 18562 20335 18590
rect 20195 18556 20335 18562
rect 20195 18528 20301 18556
rect 20229 18522 20301 18528
rect 20229 18494 20335 18522
rect 20195 18488 20335 18494
rect 20195 18460 20301 18488
rect 20229 18454 20301 18460
rect 20229 18426 20335 18454
rect 20195 18420 20335 18426
rect 20195 18392 20301 18420
rect 20229 18386 20301 18392
rect 20229 18358 20335 18386
rect 20195 18352 20335 18358
rect 20195 18324 20301 18352
rect 20229 18318 20301 18324
rect 20229 18290 20335 18318
rect 20195 18284 20335 18290
rect 20195 18256 20301 18284
rect 20229 18250 20301 18256
rect 20229 18222 20335 18250
rect 20195 18216 20335 18222
rect 20195 18188 20301 18216
rect 20229 18182 20301 18188
rect 20229 18154 20335 18182
rect 20195 18148 20335 18154
rect 20195 18120 20301 18148
rect 20229 18114 20301 18120
rect 20229 18086 20335 18114
rect 20195 18080 20335 18086
rect 20195 18052 20301 18080
rect 20229 18046 20301 18052
rect 20229 18018 20335 18046
rect 20195 18012 20335 18018
rect 20195 17984 20301 18012
rect 20229 17978 20301 17984
rect 20229 17950 20335 17978
rect 20195 17944 20335 17950
rect 20195 17916 20301 17944
rect 20229 17910 20301 17916
rect 20229 17882 20335 17910
rect 20195 17876 20335 17882
rect 20195 17848 20301 17876
rect 20229 17842 20301 17848
rect 20229 17814 20335 17842
rect 20195 17808 20335 17814
rect 20195 17780 20301 17808
rect 20229 17774 20301 17780
rect 20229 17746 20335 17774
rect 20195 17740 20335 17746
rect 20195 17712 20301 17740
rect 11457 17602 11491 17636
rect 11457 17534 11491 17568
rect 11589 17554 11623 17660
rect 12245 17554 12279 17660
rect 12351 17554 12385 17660
rect 13007 17554 13041 17660
rect 13663 17552 13697 17685
rect 14319 17552 14353 17692
rect 14975 17552 15009 17694
rect 15631 17554 15665 17681
rect 16287 17554 16321 17679
rect 17181 17672 17321 17706
rect 16393 17554 16427 17660
rect 17049 17554 17083 17660
rect 17215 17638 17287 17672
rect 17181 17604 17321 17638
rect 17215 17570 17287 17604
rect 11457 17466 11491 17500
rect 11457 17398 11491 17432
rect 11457 17330 11491 17364
rect 11457 17262 11491 17296
rect 11457 17194 11491 17228
rect 11457 17126 11491 17160
rect 11457 17058 11491 17092
rect 11457 16990 11491 17024
rect 11457 16922 11491 16956
rect 11457 16854 11491 16888
rect 11457 16786 11491 16820
rect 11457 16718 11491 16752
rect 11457 16650 11491 16684
rect 11457 16582 11491 16616
rect 11457 16514 11491 16548
rect 11457 16446 11491 16480
rect 11457 16378 11491 16412
rect 8964 16312 8988 16346
rect 9022 16312 9056 16346
rect 9090 16312 9124 16346
rect 9158 16312 9192 16346
rect 9226 16312 9260 16346
rect 9294 16312 9328 16346
rect 9362 16312 9396 16346
rect 9430 16312 9464 16346
rect 9498 16312 9532 16346
rect 9566 16312 9600 16346
rect 9634 16312 9668 16346
rect 9702 16312 9736 16346
rect 9770 16312 9804 16346
rect 9838 16322 9938 16346
rect 9838 16312 9904 16322
rect 8964 16266 8998 16312
rect 8964 16198 8998 16232
rect 9904 16254 9938 16288
rect 9791 16220 9904 16221
rect 8964 16130 8998 16164
rect 8964 16062 8998 16096
rect 9464 16186 9938 16220
rect 9464 16152 9904 16186
rect 9464 16131 9938 16152
rect 9464 16130 9814 16131
rect 9464 16033 9574 16130
rect 9704 16033 9814 16130
rect 9904 16118 9938 16131
rect 9904 16050 9938 16084
rect 8964 15994 8998 16028
rect 8964 15926 8998 15960
rect 8964 15858 8998 15892
rect 8964 15790 8998 15824
rect 8964 15722 8998 15756
rect 8964 15654 8998 15688
rect 8964 15515 8998 15620
rect 8964 15447 8998 15481
rect 8964 15379 8998 15413
rect 8964 15311 8998 15345
rect 8964 15243 8998 15277
rect 11457 16310 11491 16344
rect 11457 16242 11491 16276
rect 11457 16174 11491 16208
rect 11457 16106 11491 16140
rect 17181 17536 17321 17570
rect 17429 17554 17463 17642
rect 18085 17556 18119 17642
rect 18741 17554 18775 17708
rect 20229 17706 20301 17712
rect 20229 17678 20335 17706
rect 20195 17672 20335 17678
rect 25833 18962 25867 18996
rect 25833 18894 25867 18928
rect 25833 18826 25867 18860
rect 25833 18758 25867 18792
rect 25833 18690 25867 18724
rect 25833 18622 25867 18656
rect 25833 18554 25867 18588
rect 25833 18486 25867 18520
rect 25833 18418 25867 18452
rect 25833 18350 25867 18384
rect 25833 18282 25867 18316
rect 25833 18214 25867 18248
rect 25833 18146 25867 18180
rect 25833 18078 25867 18112
rect 25833 18010 25867 18044
rect 25833 17942 25867 17976
rect 25833 17874 25867 17908
rect 25833 17806 25867 17840
rect 25833 17738 25867 17772
rect 19397 17554 19431 17651
rect 20053 17554 20087 17651
rect 20195 17638 20301 17672
rect 20195 17604 20335 17638
rect 20195 17602 20301 17604
rect 20229 17570 20301 17602
rect 20443 17588 20477 17676
rect 21099 17588 21133 17676
rect 21755 17588 21789 17676
rect 22411 17588 22445 17676
rect 23067 17588 23101 17674
rect 23723 17588 23757 17676
rect 24379 17588 24413 17663
rect 25035 17588 25069 17676
rect 25691 17588 25725 17674
rect 25833 17670 25867 17704
rect 25833 17602 25867 17636
rect 20229 17568 20335 17570
rect 17215 17502 17287 17536
rect 17181 17468 17321 17502
rect 17215 17434 17287 17468
rect 17181 17400 17321 17434
rect 17215 17366 17287 17400
rect 17181 17332 17321 17366
rect 17215 17298 17287 17332
rect 17181 17264 17321 17298
rect 17215 17230 17287 17264
rect 17181 17196 17321 17230
rect 17215 17162 17287 17196
rect 17181 17128 17321 17162
rect 17215 17094 17287 17128
rect 17181 17060 17321 17094
rect 17215 17026 17287 17060
rect 17181 16992 17321 17026
rect 17215 16958 17287 16992
rect 17181 16924 17321 16958
rect 17215 16890 17287 16924
rect 17181 16856 17321 16890
rect 17215 16822 17287 16856
rect 17181 16788 17321 16822
rect 17215 16754 17287 16788
rect 17181 16720 17321 16754
rect 17215 16686 17287 16720
rect 17181 16652 17321 16686
rect 17215 16618 17287 16652
rect 17181 16584 17321 16618
rect 17215 16550 17287 16584
rect 17181 16516 17321 16550
rect 17215 16482 17287 16516
rect 20195 17536 20335 17568
rect 20195 17534 20301 17536
rect 20229 17502 20301 17534
rect 20229 17500 20335 17502
rect 20195 17468 20335 17500
rect 20195 17466 20301 17468
rect 20229 17434 20301 17466
rect 20229 17432 20335 17434
rect 20195 17400 20335 17432
rect 20195 17398 20301 17400
rect 20229 17366 20301 17398
rect 20229 17364 20335 17366
rect 20195 17332 20335 17364
rect 20195 17330 20301 17332
rect 20229 17298 20301 17330
rect 20229 17296 20335 17298
rect 20195 17264 20335 17296
rect 20195 17262 20301 17264
rect 20229 17230 20301 17262
rect 20229 17228 20335 17230
rect 20195 17196 20335 17228
rect 20195 17194 20301 17196
rect 20229 17162 20301 17194
rect 20229 17160 20335 17162
rect 20195 17128 20335 17160
rect 20195 17126 20301 17128
rect 20229 17094 20301 17126
rect 20229 17092 20335 17094
rect 20195 17060 20335 17092
rect 20195 17058 20301 17060
rect 20229 17026 20301 17058
rect 20229 17024 20335 17026
rect 20195 16992 20335 17024
rect 20195 16990 20301 16992
rect 20229 16958 20301 16990
rect 20229 16956 20335 16958
rect 20195 16924 20335 16956
rect 20195 16922 20301 16924
rect 20229 16890 20301 16922
rect 20229 16888 20335 16890
rect 20195 16856 20335 16888
rect 20195 16854 20301 16856
rect 20229 16822 20301 16854
rect 20229 16820 20335 16822
rect 20195 16788 20335 16820
rect 20195 16786 20301 16788
rect 20229 16754 20301 16786
rect 25833 17534 25867 17568
rect 25833 17466 25867 17500
rect 25833 17398 25867 17432
rect 25833 17330 25867 17364
rect 25833 17262 25867 17296
rect 25833 17194 25867 17228
rect 25833 17126 25867 17160
rect 25833 17058 25867 17092
rect 25833 16990 25867 17024
rect 25833 16922 25867 16956
rect 25833 16854 25867 16888
rect 25833 16786 25867 16820
rect 20229 16752 20335 16754
rect 20195 16720 20335 16752
rect 20195 16718 20301 16720
rect 20229 16686 20301 16718
rect 20229 16684 20335 16686
rect 20195 16652 20335 16684
rect 20195 16650 20301 16652
rect 20229 16618 20301 16650
rect 20229 16616 20335 16618
rect 20195 16584 20335 16616
rect 25691 16585 25725 16768
rect 25833 16718 25867 16752
rect 25833 16650 25867 16684
rect 20195 16582 20301 16584
rect 20229 16550 20301 16582
rect 20229 16548 20335 16550
rect 20195 16516 20335 16548
rect 20195 16514 20301 16516
rect 17181 16448 17321 16482
rect 17215 16414 17287 16448
rect 17181 16380 17321 16414
rect 17215 16346 17287 16380
rect 17181 16312 17321 16346
rect 17215 16278 17287 16312
rect 20053 16293 20087 16504
rect 20229 16482 20301 16514
rect 20229 16480 20335 16482
rect 20195 16448 20335 16480
rect 20195 16446 20301 16448
rect 20229 16414 20301 16446
rect 20229 16412 20335 16414
rect 20195 16380 20335 16412
rect 20195 16378 20301 16380
rect 20229 16346 20301 16378
rect 20229 16344 20335 16346
rect 20195 16312 20335 16344
rect 20195 16310 20301 16312
rect 17181 16244 17321 16278
rect 17215 16210 17287 16244
rect 17181 16176 17321 16210
rect 17215 16142 17287 16176
rect 17181 16082 17321 16142
rect 20229 16278 20301 16310
rect 20229 16276 20335 16278
rect 20195 16244 20335 16276
rect 20195 16242 20301 16244
rect 20229 16210 20301 16242
rect 25833 16582 25867 16616
rect 25833 16514 25867 16548
rect 25833 16446 25867 16480
rect 25833 16378 25867 16412
rect 25833 16310 25867 16344
rect 25833 16242 25867 16276
rect 20229 16208 20335 16210
rect 20195 16176 20335 16208
rect 24379 16196 24413 16238
rect 20195 16174 20301 16176
rect 20229 16142 20301 16174
rect 24368 16150 24424 16196
rect 25833 16174 25867 16208
rect 20229 16140 20335 16142
rect 20195 16106 20335 16140
rect 11491 16072 11581 16082
rect 11457 16048 11581 16072
rect 11615 16048 11649 16082
rect 11683 16048 11717 16082
rect 11751 16048 11785 16082
rect 11819 16048 11853 16082
rect 11887 16048 11921 16082
rect 11955 16048 11989 16082
rect 12023 16048 12057 16082
rect 12091 16048 12125 16082
rect 12159 16048 12193 16082
rect 12227 16048 12261 16082
rect 12295 16048 12329 16082
rect 12363 16048 12397 16082
rect 12431 16048 12465 16082
rect 12499 16048 12533 16082
rect 12567 16048 12601 16082
rect 12635 16048 12669 16082
rect 12703 16048 12737 16082
rect 12771 16048 12805 16082
rect 12839 16048 12873 16082
rect 12907 16048 12941 16082
rect 12975 16048 13009 16082
rect 13043 16048 13077 16082
rect 13111 16048 13145 16082
rect 13179 16048 13213 16082
rect 13247 16048 13281 16082
rect 13315 16048 13349 16082
rect 13383 16048 13417 16082
rect 13451 16048 13485 16082
rect 13519 16048 13553 16082
rect 13587 16048 13621 16082
rect 13655 16048 13689 16082
rect 13723 16048 13757 16082
rect 13791 16048 13825 16082
rect 13859 16048 13893 16082
rect 13927 16048 13961 16082
rect 13995 16048 14029 16082
rect 14063 16048 14097 16082
rect 14131 16048 14165 16082
rect 14199 16048 14233 16082
rect 14267 16048 14301 16082
rect 14335 16048 14369 16082
rect 14403 16048 14437 16082
rect 14471 16048 14505 16082
rect 14539 16048 14573 16082
rect 14607 16048 14641 16082
rect 14675 16048 14709 16082
rect 14743 16048 14777 16082
rect 14811 16048 14845 16082
rect 14879 16048 14913 16082
rect 14947 16048 14981 16082
rect 15015 16048 15049 16082
rect 15083 16048 15117 16082
rect 15151 16048 15185 16082
rect 15219 16048 15253 16082
rect 15287 16048 15321 16082
rect 15355 16048 15389 16082
rect 15423 16048 15457 16082
rect 15491 16048 15525 16082
rect 15559 16048 15593 16082
rect 15627 16048 15661 16082
rect 15695 16048 15729 16082
rect 15763 16048 15797 16082
rect 15831 16048 15865 16082
rect 15899 16048 15933 16082
rect 15967 16048 16001 16082
rect 16035 16048 16069 16082
rect 16103 16048 16137 16082
rect 16171 16048 16205 16082
rect 16239 16048 16273 16082
rect 16307 16048 16341 16082
rect 16375 16048 16409 16082
rect 16443 16048 16477 16082
rect 16511 16048 16545 16082
rect 16579 16048 16613 16082
rect 16647 16048 16681 16082
rect 16715 16048 16749 16082
rect 16783 16048 16817 16082
rect 16851 16048 16885 16082
rect 16919 16048 16953 16082
rect 16987 16048 17021 16082
rect 17055 16048 17089 16082
rect 17123 16048 17157 16082
rect 17191 16048 17311 16082
rect 17345 16048 17379 16082
rect 17413 16048 17447 16082
rect 17481 16048 17515 16082
rect 17549 16048 17583 16082
rect 17617 16048 17651 16082
rect 17685 16048 17719 16082
rect 17753 16048 17787 16082
rect 17821 16048 17855 16082
rect 17889 16048 17923 16082
rect 17957 16048 17991 16082
rect 18025 16048 18059 16082
rect 18093 16048 18127 16082
rect 18161 16048 18195 16082
rect 18229 16048 18263 16082
rect 18297 16048 18331 16082
rect 18365 16048 18399 16082
rect 18433 16048 18467 16082
rect 18501 16048 18535 16082
rect 18569 16048 18603 16082
rect 18637 16048 18671 16082
rect 18705 16048 18739 16082
rect 18773 16048 18807 16082
rect 18841 16048 18875 16082
rect 18909 16048 18943 16082
rect 18977 16048 19011 16082
rect 19045 16048 19079 16082
rect 19113 16048 19147 16082
rect 19181 16048 19215 16082
rect 19249 16048 19283 16082
rect 19317 16048 19351 16082
rect 19385 16048 19419 16082
rect 19453 16048 19487 16082
rect 19521 16048 19555 16082
rect 19589 16048 19623 16082
rect 19657 16048 19691 16082
rect 19725 16048 19759 16082
rect 19793 16048 19827 16082
rect 19861 16048 19895 16082
rect 19929 16048 19963 16082
rect 19997 16048 20031 16082
rect 20065 16048 20099 16082
rect 20133 16072 20195 16082
rect 20229 16082 20335 16106
rect 25833 16106 25867 16140
rect 20229 16072 20325 16082
rect 20133 16048 20325 16072
rect 20359 16048 20393 16082
rect 20427 16048 20461 16082
rect 20495 16048 20529 16082
rect 20563 16048 20597 16082
rect 20631 16048 20665 16082
rect 20699 16048 20733 16082
rect 20767 16048 20801 16082
rect 20835 16048 20869 16082
rect 20903 16048 20937 16082
rect 20971 16048 21005 16082
rect 21039 16048 21073 16082
rect 21107 16048 21141 16082
rect 21175 16048 21209 16082
rect 21243 16048 21277 16082
rect 21311 16048 21345 16082
rect 21379 16048 21413 16082
rect 21447 16048 21481 16082
rect 21515 16048 21549 16082
rect 21583 16048 21617 16082
rect 21651 16048 21685 16082
rect 21719 16048 21753 16082
rect 21787 16048 21821 16082
rect 21855 16048 21889 16082
rect 21923 16048 21957 16082
rect 21991 16048 22025 16082
rect 22059 16048 22093 16082
rect 22127 16048 22161 16082
rect 22195 16048 22229 16082
rect 22263 16048 22297 16082
rect 22331 16048 22365 16082
rect 22399 16048 22433 16082
rect 22467 16048 22501 16082
rect 22535 16048 22569 16082
rect 22603 16048 22637 16082
rect 22671 16048 22705 16082
rect 22739 16048 22773 16082
rect 22807 16048 22841 16082
rect 22875 16048 22909 16082
rect 22943 16048 22977 16082
rect 23011 16048 23045 16082
rect 23079 16048 23113 16082
rect 23147 16048 23181 16082
rect 23215 16048 23249 16082
rect 23283 16048 23317 16082
rect 23351 16048 23385 16082
rect 23419 16048 23453 16082
rect 23487 16048 23521 16082
rect 23555 16048 23589 16082
rect 23623 16048 23657 16082
rect 23691 16048 23725 16082
rect 23759 16048 23793 16082
rect 23827 16048 23861 16082
rect 23895 16048 23929 16082
rect 23963 16048 23997 16082
rect 24031 16048 24065 16082
rect 24099 16048 24133 16082
rect 24167 16048 24201 16082
rect 24235 16048 24269 16082
rect 24303 16048 24337 16082
rect 24371 16048 24405 16082
rect 24439 16048 24473 16082
rect 24507 16048 24541 16082
rect 24575 16048 24609 16082
rect 24643 16048 24677 16082
rect 24711 16048 24745 16082
rect 24779 16048 24813 16082
rect 24847 16048 24881 16082
rect 24915 16048 24949 16082
rect 24983 16048 25017 16082
rect 25051 16048 25085 16082
rect 25119 16048 25153 16082
rect 25187 16048 25221 16082
rect 25255 16048 25289 16082
rect 25323 16048 25357 16082
rect 25391 16048 25425 16082
rect 25459 16048 25493 16082
rect 25527 16048 25561 16082
rect 25595 16048 25629 16082
rect 25663 16048 25697 16082
rect 25731 16048 25765 16082
rect 25799 16072 25833 16082
rect 25799 16048 25867 16072
rect 9904 15982 9938 16016
rect 11458 15976 11516 16048
rect 13704 15976 13762 16048
rect 9904 15914 9938 15948
rect 9904 15846 9938 15880
rect 9904 15778 9938 15812
rect 9904 15710 9938 15744
rect 9904 15642 9938 15676
rect 9904 15574 9938 15608
rect 9904 15506 9938 15540
rect 9904 15438 9938 15472
rect 9904 15370 9938 15404
rect 9904 15302 9938 15336
rect 11457 15942 11481 15976
rect 11515 15942 11549 15976
rect 11583 15942 11617 15976
rect 11651 15942 11685 15976
rect 11719 15942 11753 15976
rect 11787 15942 11821 15976
rect 11855 15942 11889 15976
rect 11923 15942 11957 15976
rect 11991 15942 12025 15976
rect 12059 15942 12093 15976
rect 12127 15942 12161 15976
rect 12195 15942 12229 15976
rect 12263 15942 12297 15976
rect 12331 15942 12365 15976
rect 12399 15942 12433 15976
rect 12467 15942 12501 15976
rect 12535 15942 12649 15976
rect 12683 15942 12717 15976
rect 12751 15942 12785 15976
rect 12819 15942 12853 15976
rect 12887 15942 12921 15976
rect 12955 15942 12989 15976
rect 13023 15942 13057 15976
rect 13091 15942 13125 15976
rect 13159 15942 13193 15976
rect 13227 15942 13261 15976
rect 13295 15942 13329 15976
rect 13363 15942 13397 15976
rect 13431 15942 13465 15976
rect 13499 15942 13533 15976
rect 13567 15942 13601 15976
rect 13635 15942 13669 15976
rect 13703 15952 13793 15976
rect 13866 15974 13924 16048
rect 14862 15974 14932 16048
rect 15004 15975 15074 16048
rect 18112 15976 18204 16048
rect 17215 15975 17239 15976
rect 13703 15942 13759 15952
rect 11457 15902 11491 15942
rect 11457 15834 11491 15868
rect 13759 15884 13793 15918
rect 13759 15816 13793 15850
rect 13386 15811 13759 15812
rect 11457 15766 11491 15800
rect 11457 15722 11491 15732
rect 11787 15765 11853 15811
rect 12018 15765 12134 15811
rect 12265 15765 12333 15811
rect 11787 15723 11821 15765
rect 11457 15698 11710 15722
rect 12043 15712 12077 15765
rect 12299 15723 12333 15765
rect 12917 15765 13006 15811
rect 13129 15765 13264 15811
rect 13375 15782 13759 15811
rect 13375 15765 13793 15782
rect 12917 15704 12951 15765
rect 11491 15664 11710 15698
rect 13173 15695 13207 15765
rect 13386 15764 13793 15765
rect 13429 15723 13463 15764
rect 13759 15748 13793 15764
rect 11457 15630 11710 15664
rect 11491 15596 11710 15630
rect 13759 15680 13793 15714
rect 13759 15612 13793 15646
rect 11457 15562 11491 15596
rect 11457 15494 11491 15528
rect 11457 15426 11491 15460
rect 11457 15358 11491 15392
rect 11457 15290 11491 15324
rect 10595 15268 10671 15287
rect 9904 15234 9938 15268
rect 8998 15209 9354 15216
rect 8964 15175 9354 15209
rect 8998 15160 9354 15175
rect 8964 15107 8998 15141
rect 9154 15097 9354 15160
rect 9904 15166 9938 15200
rect 9904 15098 9938 15132
rect 8964 15039 8998 15073
rect 9616 15011 9662 15038
rect 9904 15030 9938 15064
rect 8964 14971 8998 15005
rect 9354 14977 9662 15011
rect 9704 14977 9814 15011
rect 8964 14903 8998 14937
rect 9904 14962 9938 14996
rect 10046 15258 10450 15268
rect 10046 15224 10329 15258
rect 10363 15224 10450 15258
rect 10046 15208 10450 15224
rect 10595 15234 10618 15268
rect 10652 15234 10671 15268
rect 10595 15215 10671 15234
rect 13759 15544 13793 15578
rect 13759 15476 13793 15510
rect 13759 15408 13793 15442
rect 13759 15340 13793 15374
rect 11457 15222 11491 15256
rect 10046 15012 10106 15208
rect 10257 15117 10312 15171
rect 10260 15030 10294 15117
rect 10468 15024 10502 15170
rect 10676 15042 10710 15120
rect 10741 15117 10796 15171
rect 10956 15027 10990 15167
rect 11457 15154 11491 15188
rect 11457 15086 11491 15120
rect 10046 14978 10057 15012
rect 10091 14978 10106 15012
rect 10046 14964 10106 14978
rect 11457 15018 11491 15052
rect 11787 15081 11821 15136
rect 12043 15081 12077 15136
rect 12555 15081 12589 15286
rect 13759 15272 13793 15306
rect 13759 15204 13793 15238
rect 13429 15081 13463 15141
rect 11787 15035 11900 15081
rect 12003 15035 12088 15081
rect 12515 15035 12589 15081
rect 13352 15035 13463 15081
rect 13759 15136 13793 15170
rect 13759 15068 13793 15102
rect 9904 14879 9938 14928
rect 11457 14950 11491 14984
rect 11457 14882 11491 14916
rect 8998 14869 9064 14879
rect 8964 14845 9064 14869
rect 9098 14845 9132 14879
rect 9166 14845 9200 14879
rect 9234 14845 9268 14879
rect 9302 14845 9336 14879
rect 9370 14845 9404 14879
rect 9438 14845 9472 14879
rect 9506 14845 9540 14879
rect 9574 14845 9608 14879
rect 9642 14845 9676 14879
rect 9710 14845 9744 14879
rect 9778 14845 9812 14879
rect 9846 14845 9880 14879
rect 9914 14845 9938 14879
rect 9526 14800 9574 14802
rect 10086 14800 10134 14818
rect 9526 14796 10134 14800
rect 9526 14762 9533 14796
rect 9567 14795 10134 14796
rect 9567 14762 10090 14795
rect 9526 14761 10090 14762
rect 10124 14761 10134 14795
rect 10174 14807 10208 14847
rect 10346 14810 10380 14847
rect 10346 14807 10518 14810
rect 10174 14796 10518 14807
rect 10174 14773 10458 14796
rect 9526 14756 10134 14761
rect 9526 14754 9574 14756
rect 10086 14740 10134 14756
rect 10346 14762 10458 14773
rect 10492 14762 10518 14796
rect 10346 14750 10518 14762
rect 9650 14716 9674 14722
rect 8964 14682 8988 14716
rect 9022 14682 9056 14716
rect 9090 14682 9124 14716
rect 9158 14682 9192 14716
rect 9226 14682 9260 14716
rect 9294 14682 9328 14716
rect 9362 14682 9396 14716
rect 9430 14682 9464 14716
rect 9498 14682 9532 14716
rect 9566 14688 9674 14716
rect 9708 14688 9742 14722
rect 9776 14688 9810 14722
rect 9844 14716 9936 14722
rect 9844 14688 9926 14716
rect 9566 14682 9684 14688
rect 9902 14682 9926 14688
rect 9960 14682 10048 14716
rect 10346 14715 10380 14750
rect 8964 14600 8998 14682
rect 10014 14664 10048 14682
rect 10332 14681 10380 14715
rect 10554 14681 10588 14862
rect 10834 14810 10868 14865
rect 10834 14798 11000 14810
rect 10748 14794 11000 14798
rect 10748 14760 10938 14794
rect 10972 14760 11000 14794
rect 10748 14750 11000 14760
rect 11041 14808 11075 14881
rect 13759 15000 13793 15034
rect 13759 14932 13793 14966
rect 13759 14858 13793 14898
rect 11491 14848 11559 14858
rect 11457 14824 11559 14848
rect 11593 14824 11627 14858
rect 11661 14824 11695 14858
rect 11729 14824 11763 14858
rect 11797 14824 11831 14858
rect 11865 14824 11899 14858
rect 11933 14824 11967 14858
rect 12001 14824 12035 14858
rect 12069 14824 12103 14858
rect 12137 14824 12171 14858
rect 12205 14824 12239 14858
rect 12273 14824 12307 14858
rect 12341 14824 12375 14858
rect 12409 14824 12443 14858
rect 12477 14824 12511 14858
rect 12545 14824 12579 14858
rect 12613 14824 12647 14858
rect 12681 14824 12715 14858
rect 12749 14824 12783 14858
rect 12817 14824 12851 14858
rect 12885 14824 12919 14858
rect 12953 14824 12987 14858
rect 13021 14824 13055 14858
rect 13089 14824 13123 14858
rect 13157 14824 13191 14858
rect 13225 14824 13259 14858
rect 13293 14824 13327 14858
rect 13361 14824 13395 14858
rect 13429 14824 13463 14858
rect 13497 14824 13531 14858
rect 13565 14824 13599 14858
rect 13633 14824 13667 14858
rect 13701 14824 13735 14858
rect 13769 14824 13793 14858
rect 13865 15940 13889 15974
rect 13923 15940 13957 15974
rect 13991 15940 14025 15974
rect 14059 15940 14093 15974
rect 14127 15940 14161 15974
rect 14195 15940 14229 15974
rect 14263 15940 14297 15974
rect 14331 15940 14365 15974
rect 14399 15940 14433 15974
rect 14467 15940 14501 15974
rect 14535 15940 14569 15974
rect 14603 15940 14637 15974
rect 14671 15940 14705 15974
rect 14739 15940 14773 15974
rect 14807 15958 14932 15974
rect 14807 15950 14931 15958
rect 14807 15940 14897 15950
rect 13865 15872 13899 15940
rect 14897 15882 14931 15916
rect 13865 15865 13988 15872
rect 13899 15861 13988 15865
rect 13899 15831 14009 15861
rect 13865 15818 14009 15831
rect 14208 15818 14549 15872
rect 14778 15848 14897 15872
rect 15003 15941 15027 15975
rect 15061 15941 15095 15975
rect 15129 15941 15163 15975
rect 15197 15941 15231 15975
rect 15265 15941 15299 15975
rect 15333 15941 15367 15975
rect 15401 15941 15435 15975
rect 15469 15941 15503 15975
rect 15537 15941 15571 15975
rect 15605 15941 15639 15975
rect 15673 15941 15707 15975
rect 15741 15941 15775 15975
rect 15809 15941 15843 15975
rect 15877 15941 15911 15975
rect 15945 15941 15979 15975
rect 16013 15941 16047 15975
rect 16081 15941 16115 15975
rect 16149 15941 16183 15975
rect 16217 15941 16251 15975
rect 16285 15941 16319 15975
rect 16353 15941 16387 15975
rect 16421 15941 16455 15975
rect 16489 15941 16523 15975
rect 16557 15941 16591 15975
rect 16625 15941 16659 15975
rect 16693 15941 16727 15975
rect 16761 15941 16795 15975
rect 16829 15941 16863 15975
rect 16897 15941 16931 15975
rect 16965 15941 16999 15975
rect 17033 15941 17067 15975
rect 17101 15941 17135 15975
rect 17169 15942 17239 15975
rect 17273 15942 17307 15976
rect 17341 15942 17375 15976
rect 17409 15942 17443 15976
rect 17477 15942 17511 15976
rect 17545 15942 17579 15976
rect 17613 15942 17647 15976
rect 17681 15942 17715 15976
rect 17749 15942 17783 15976
rect 17817 15942 17851 15976
rect 17885 15942 17919 15976
rect 17953 15942 17987 15976
rect 18021 15942 18055 15976
rect 18089 15952 18205 15976
rect 18089 15942 18171 15952
rect 17169 15941 17249 15942
rect 15003 15902 15037 15941
rect 14931 15868 15003 15872
rect 18171 15884 18205 15918
rect 15037 15868 15038 15872
rect 14931 15854 15038 15868
rect 14931 15848 17793 15854
rect 14778 15834 17793 15848
rect 14778 15818 15003 15834
rect 13865 15797 13899 15818
rect 13865 15729 13899 15763
rect 13975 15716 14009 15818
rect 14487 15725 14521 15818
rect 14886 15814 15003 15818
rect 14886 15800 14897 15814
rect 14931 15800 15003 15814
rect 15037 15800 17793 15834
rect 17892 15850 18171 15854
rect 17892 15816 18205 15850
rect 17892 15800 18171 15816
rect 14897 15746 14931 15780
rect 13865 15661 13899 15695
rect 13865 15593 13899 15627
rect 13865 15525 13899 15559
rect 13865 15457 13899 15491
rect 13865 15358 13899 15423
rect 13865 15290 13899 15324
rect 13865 15222 13899 15256
rect 13865 15154 13899 15188
rect 13865 15086 13899 15120
rect 13865 15018 13899 15052
rect 13865 14950 13899 14984
rect 13865 14882 13899 14916
rect 14897 15678 14931 15712
rect 14897 15610 14931 15644
rect 14897 15542 14931 15576
rect 14897 15474 14931 15508
rect 14897 15406 14931 15440
rect 14897 15338 14931 15372
rect 14897 15270 14931 15304
rect 14897 15202 14931 15236
rect 14897 15134 14931 15168
rect 14897 15066 14931 15100
rect 14897 14998 14931 15032
rect 14897 14930 14931 14964
rect 14897 14858 14931 14896
rect 13899 14848 13989 14858
rect 13865 14824 13989 14848
rect 14023 14824 14057 14858
rect 14091 14824 14125 14858
rect 14159 14824 14193 14858
rect 14227 14824 14261 14858
rect 14295 14824 14329 14858
rect 14363 14824 14397 14858
rect 14431 14824 14465 14858
rect 14499 14824 14533 14858
rect 14567 14824 14601 14858
rect 14635 14824 14669 14858
rect 14703 14824 14737 14858
rect 14771 14824 14805 14858
rect 14839 14824 14873 14858
rect 14907 14824 14931 14858
rect 15003 15766 15037 15800
rect 15003 15698 15037 15732
rect 15109 15704 15143 15800
rect 15765 15730 15799 15800
rect 16543 15695 16577 15800
rect 17321 15730 17355 15800
rect 17977 15730 18011 15800
rect 18171 15748 18205 15782
rect 15003 15630 15037 15664
rect 15003 15562 15037 15596
rect 18171 15680 18205 15714
rect 18171 15612 18205 15646
rect 21241 15617 21352 15817
rect 21404 15617 21438 15817
rect 15003 15494 15037 15528
rect 15887 15471 15921 15577
rect 18171 15544 18205 15578
rect 18171 15476 18205 15510
rect 15003 15426 15037 15460
rect 15003 15358 15037 15392
rect 15003 15290 15037 15324
rect 15003 15222 15037 15256
rect 15003 15154 15037 15188
rect 15003 15086 15037 15120
rect 21342 15506 21412 15526
rect 21342 15472 21360 15506
rect 21394 15472 21412 15506
rect 21342 15454 21412 15472
rect 18171 15408 18205 15442
rect 18171 15340 18205 15374
rect 18171 15272 18205 15306
rect 18171 15204 18205 15238
rect 18171 15136 18205 15170
rect 18171 15068 18205 15102
rect 15003 15018 15037 15052
rect 15003 14950 15037 14984
rect 15109 15013 15143 15055
rect 15765 15013 15799 15055
rect 17199 15013 17233 15055
rect 15109 14967 15228 15013
rect 15693 14967 15799 15013
rect 17169 14967 17233 15013
rect 17321 15013 17355 15055
rect 17977 15013 18011 15055
rect 17321 14967 17441 15013
rect 17931 14967 18011 15013
rect 18171 15000 18205 15034
rect 15003 14882 15037 14916
rect 18171 14932 18205 14966
rect 18171 14858 18205 14898
rect 15037 14848 15118 14858
rect 15003 14824 15118 14848
rect 15152 14824 15186 14858
rect 15220 14824 15254 14858
rect 15288 14824 15322 14858
rect 15356 14824 15390 14858
rect 15424 14824 15458 14858
rect 15492 14824 15526 14858
rect 15560 14824 15594 14858
rect 15628 14824 15662 14858
rect 15696 14824 15730 14858
rect 15764 14824 15798 14858
rect 15832 14824 15866 14858
rect 15900 14824 15934 14858
rect 15968 14824 16002 14858
rect 16036 14824 16070 14858
rect 16104 14824 16138 14858
rect 16172 14824 16206 14858
rect 16240 14824 16274 14858
rect 16308 14824 16342 14858
rect 16376 14824 16410 14858
rect 16444 14824 16478 14858
rect 16512 14824 16546 14858
rect 16580 14824 16651 14858
rect 16685 14824 16719 14858
rect 16753 14824 16787 14858
rect 16821 14824 16855 14858
rect 16889 14824 16923 14858
rect 16957 14824 16991 14858
rect 17025 14824 17059 14858
rect 17093 14824 17127 14858
rect 17161 14824 17195 14858
rect 17229 14824 17263 14858
rect 17297 14824 17331 14858
rect 17365 14824 17399 14858
rect 17433 14824 17467 14858
rect 17501 14824 17535 14858
rect 17569 14824 17603 14858
rect 17637 14824 17671 14858
rect 17705 14824 17739 14858
rect 17773 14824 17807 14858
rect 17841 14824 17875 14858
rect 17909 14824 17943 14858
rect 17977 14824 18011 14858
rect 18045 14824 18079 14858
rect 18113 14824 18147 14858
rect 18181 14824 18205 14858
rect 11041 14794 11158 14808
rect 11041 14760 11108 14794
rect 11142 14760 11158 14794
rect 10748 14715 10782 14750
rect 11041 14744 11158 14760
rect 11041 14682 11075 14744
rect 9378 14617 9458 14648
rect 10014 14640 10084 14664
rect 10014 14630 10050 14640
rect 8964 14532 8998 14566
rect 9154 14558 9254 14592
rect 9378 14583 9401 14617
rect 9435 14583 9458 14617
rect 9378 14558 9458 14583
rect 9582 14594 9960 14628
rect 9582 14527 9616 14594
rect 9754 14532 9788 14594
rect 9926 14539 9960 14594
rect 10050 14572 10084 14606
rect 11446 14628 11470 14662
rect 11504 14628 11538 14662
rect 11572 14628 11606 14662
rect 11640 14628 11674 14662
rect 11708 14628 11742 14662
rect 11776 14628 11810 14662
rect 11844 14628 11878 14662
rect 11912 14628 11946 14662
rect 11980 14628 12014 14662
rect 12048 14628 12082 14662
rect 12116 14628 12150 14662
rect 12184 14628 12218 14662
rect 12252 14628 12286 14662
rect 12320 14628 12354 14662
rect 12388 14628 12422 14662
rect 12456 14628 12490 14662
rect 12524 14628 12558 14662
rect 12592 14628 12626 14662
rect 12660 14628 12694 14662
rect 12728 14628 12762 14662
rect 12796 14628 12830 14662
rect 12864 14628 12898 14662
rect 12932 14628 12966 14662
rect 13000 14628 13034 14662
rect 13068 14628 13102 14662
rect 13136 14628 13170 14662
rect 13204 14638 13434 14662
rect 13204 14628 13254 14638
rect 8964 14464 8998 14498
rect 8964 14396 8998 14430
rect 8964 14328 8998 14362
rect 8964 14260 8998 14294
rect 8964 14192 8998 14226
rect 8964 14124 8998 14158
rect 8964 14056 8998 14090
rect 8964 13988 8998 14022
rect 8964 13920 8998 13954
rect 8964 13852 8998 13886
rect 8964 13784 8998 13818
rect 8964 13716 8998 13750
rect 8964 13648 8998 13682
rect 8964 13580 8998 13614
rect 8866 13522 8890 13556
rect 8924 13546 8964 13556
rect 8924 13522 8998 13546
rect 10050 14504 10084 14538
rect 10542 14570 10602 14584
rect 10542 14536 10554 14570
rect 10588 14536 10602 14570
rect 11446 14551 11480 14628
rect 10050 14446 10084 14470
rect 10174 14446 10208 14515
rect 10468 14446 10502 14522
rect 10542 14518 10602 14536
rect 10662 14446 10696 14530
rect 10834 14446 10868 14537
rect 10955 14446 10989 14539
rect 13288 14628 13342 14638
rect 13254 14570 13288 14604
rect 11480 14517 11635 14544
rect 11446 14490 11635 14517
rect 11941 14490 12843 14544
rect 13376 14628 13434 14638
rect 13468 14628 13502 14662
rect 13536 14628 13570 14662
rect 13604 14628 13638 14662
rect 13672 14628 13706 14662
rect 13740 14628 13774 14662
rect 13808 14628 13842 14662
rect 13876 14628 13910 14662
rect 13944 14628 13978 14662
rect 14012 14628 14046 14662
rect 14080 14628 14114 14662
rect 14148 14628 14182 14662
rect 14216 14628 14250 14662
rect 14284 14628 14318 14662
rect 14352 14628 14386 14662
rect 14420 14628 14454 14662
rect 14488 14628 14522 14662
rect 14556 14628 14590 14662
rect 14624 14628 14658 14662
rect 14692 14628 14726 14662
rect 14760 14628 14794 14662
rect 14828 14628 14862 14662
rect 14896 14628 14930 14662
rect 14964 14628 14998 14662
rect 15032 14628 15066 14662
rect 15100 14628 15134 14662
rect 15168 14628 15202 14662
rect 15236 14628 15270 14662
rect 15304 14628 15338 14662
rect 15372 14628 15406 14662
rect 15440 14628 15474 14662
rect 15508 14628 15542 14662
rect 15576 14628 15610 14662
rect 15644 14628 15678 14662
rect 15712 14628 15746 14662
rect 15780 14628 15814 14662
rect 15848 14628 15882 14662
rect 15916 14628 15950 14662
rect 15984 14628 16018 14662
rect 16052 14628 16086 14662
rect 16120 14628 16154 14662
rect 16188 14628 16222 14662
rect 16256 14628 16290 14662
rect 16324 14628 16358 14662
rect 16392 14628 16426 14662
rect 16460 14628 16494 14662
rect 16528 14628 16562 14662
rect 16596 14628 16630 14662
rect 16664 14628 16698 14662
rect 16732 14628 16766 14662
rect 16800 14628 16834 14662
rect 16868 14628 16902 14662
rect 16936 14628 16970 14662
rect 17004 14628 17038 14662
rect 17072 14628 17106 14662
rect 17140 14628 17174 14662
rect 17208 14628 17242 14662
rect 17276 14628 17310 14662
rect 17344 14628 17378 14662
rect 17412 14628 17446 14662
rect 17480 14628 17514 14662
rect 17548 14628 17582 14662
rect 17616 14628 17650 14662
rect 17684 14628 17718 14662
rect 17752 14628 17786 14662
rect 17820 14628 17854 14662
rect 17888 14628 17922 14662
rect 17956 14628 17990 14662
rect 18024 14628 18058 14662
rect 18092 14628 18126 14662
rect 18160 14628 18194 14662
rect 18228 14628 18262 14662
rect 18296 14628 18330 14662
rect 18364 14628 18388 14662
rect 13342 14570 13376 14604
rect 13254 14502 13288 14536
rect 13338 14536 13342 14560
rect 18354 14594 18388 14628
rect 13376 14536 13581 14560
rect 13338 14514 13581 14536
rect 15236 14514 15310 14560
rect 16330 14514 16403 14560
rect 18198 14526 18388 14560
rect 18198 14514 18354 14526
rect 11446 14483 11480 14490
rect 11446 14446 11480 14449
rect 10050 14436 11480 14446
rect 10084 14415 11480 14436
rect 10084 14402 11446 14415
rect 10050 14386 11446 14402
rect 10050 14368 10084 14386
rect 10050 14300 10084 14334
rect 10882 14334 10950 14350
rect 10882 14300 10898 14334
rect 10932 14300 10950 14334
rect 10882 14280 10950 14300
rect 11446 14347 11480 14381
rect 10050 14232 10084 14266
rect 10050 14164 10084 14198
rect 10050 14096 10084 14130
rect 10050 14028 10084 14062
rect 10050 13960 10084 13994
rect 10050 13892 10084 13926
rect 10050 13824 10084 13858
rect 10050 13756 10084 13790
rect 10050 13688 10084 13722
rect 10050 13587 10084 13654
rect 8866 13451 8900 13522
rect 10050 13519 10084 13553
rect 8866 13383 8900 13417
rect 8866 13315 8900 13349
rect 8866 13247 8900 13281
rect 9154 13223 9254 13512
rect 10050 13451 10084 13485
rect 10050 13383 10084 13417
rect 10050 13315 10084 13349
rect 10050 13247 10084 13281
rect 8900 13213 8940 13223
rect 8866 13189 8940 13213
rect 8974 13189 9008 13223
rect 9042 13189 9076 13223
rect 9110 13189 9144 13223
rect 9178 13189 9212 13223
rect 9246 13189 9280 13223
rect 9314 13189 9348 13223
rect 9382 13189 9406 13223
rect 9372 13092 9406 13189
rect 9372 13024 9406 13058
rect 9372 12956 9406 12990
rect 9372 12888 9406 12922
rect 9372 12820 9406 12854
rect 9372 12752 9406 12786
rect 9372 12684 9406 12718
rect 9372 12616 9406 12650
rect 9343 12582 9372 12592
rect 10050 13179 10084 13213
rect 10050 13111 10084 13145
rect 10050 13043 10084 13077
rect 10050 12975 10084 13009
rect 10050 12907 10084 12941
rect 10050 12839 10084 12873
rect 10050 12771 10084 12805
rect 10050 12703 10084 12737
rect 10050 12592 10084 12669
rect 11446 14279 11480 14313
rect 11446 14211 11480 14245
rect 13254 14434 13288 14468
rect 13254 14366 13288 14400
rect 13254 14298 13288 14332
rect 13254 14230 13288 14264
rect 13066 14202 13150 14214
rect 13066 14197 13103 14202
rect 13065 14184 13103 14197
rect 11446 14143 11480 14177
rect 13066 14168 13103 14184
rect 13137 14168 13150 14202
rect 13066 14154 13150 14168
rect 13254 14162 13288 14196
rect 11446 14075 11480 14109
rect 11446 14007 11480 14041
rect 11446 13939 11480 13973
rect 11446 13871 11480 13905
rect 11446 13803 11480 13837
rect 11446 13735 11480 13769
rect 11446 13667 11480 13701
rect 11446 13599 11480 13633
rect 11446 13531 11480 13565
rect 11446 13463 11480 13497
rect 11446 13395 11480 13429
rect 11446 13327 11480 13361
rect 11446 13259 11480 13293
rect 11446 13191 11480 13225
rect 11446 13123 11480 13157
rect 11446 13055 11480 13089
rect 11446 12987 11480 13021
rect 11446 12919 11480 12953
rect 11446 12818 11480 12885
rect 11446 12750 11480 12784
rect 11446 12682 11480 12716
rect 11446 12614 11480 12648
rect 9343 12558 9406 12582
rect 9343 12534 9377 12558
rect 9128 12475 9377 12534
rect 9128 12369 9191 12475
rect 9297 12474 9377 12475
rect 9496 12474 9530 12554
rect 9668 12474 9702 12585
rect 10050 12568 10113 12592
rect 10050 12558 10079 12568
rect 9840 12474 9874 12546
rect 10079 12500 10113 12534
rect 9297 12467 10079 12474
rect 9297 12433 9343 12467
rect 9377 12466 10079 12467
rect 9377 12433 10113 12466
rect 9297 12432 10113 12433
rect 9297 12420 10079 12432
rect 9297 12399 9377 12420
rect 9297 12369 9343 12399
rect 9128 12365 9343 12369
rect 9128 12331 9377 12365
rect 9128 12302 9343 12331
rect 10079 12307 10113 12398
rect 9377 12297 9443 12307
rect 9343 12273 9443 12297
rect 9477 12273 9511 12307
rect 9545 12273 9579 12307
rect 9613 12273 9647 12307
rect 9681 12273 9715 12307
rect 9749 12273 9783 12307
rect 9817 12273 9851 12307
rect 9885 12273 9919 12307
rect 9953 12273 9987 12307
rect 10021 12273 10055 12307
rect 10089 12273 10113 12307
rect 11446 12546 11480 12580
rect 11446 12478 11480 12512
rect 11446 12410 11480 12444
rect 11446 12342 11480 12376
rect 11446 12274 11480 12308
rect 11446 12206 11480 12240
rect 11446 12138 11480 12172
rect 11446 12070 11480 12104
rect 11446 12002 11480 12036
rect 11446 11934 11480 11968
rect 11446 11866 11480 11900
rect 11446 11798 11480 11832
rect 13254 14094 13288 14128
rect 13254 14026 13288 14060
rect 13254 13958 13288 13992
rect 13254 13890 13288 13924
rect 13254 13822 13288 13856
rect 13254 13754 13288 13788
rect 13254 13686 13288 13720
rect 13254 13618 13288 13652
rect 13254 13550 13288 13584
rect 13254 13482 13288 13516
rect 13254 13414 13288 13448
rect 13254 13346 13288 13380
rect 13254 13278 13288 13312
rect 13254 13210 13288 13244
rect 13342 14502 13376 14514
rect 13342 14434 13376 14468
rect 13462 14459 13496 14514
rect 15236 14447 15270 14514
rect 16348 14472 16382 14514
rect 18226 14472 18260 14514
rect 18354 14458 18388 14492
rect 13342 14366 13376 14400
rect 13342 14298 13376 14332
rect 13342 14230 13376 14264
rect 13342 14162 13376 14196
rect 13342 14094 13376 14128
rect 13342 14026 13376 14060
rect 18354 14390 18388 14424
rect 18354 14322 18388 14356
rect 18354 14254 18388 14288
rect 18354 14186 18388 14220
rect 18354 14118 18388 14152
rect 18354 14050 18388 14084
rect 13342 13958 13376 13992
rect 13342 13890 13376 13924
rect 13462 13886 13496 14004
rect 14018 13868 14052 14006
rect 14574 13907 14608 14006
rect 15130 13886 15164 13972
rect 15236 13886 15270 13972
rect 15792 13886 15826 14006
rect 16348 13889 16382 14006
rect 16452 13892 16486 13972
rect 17008 13876 17042 13972
rect 17114 13887 17148 14006
rect 18354 13982 18388 14016
rect 17670 13886 17704 13976
rect 18226 13886 18260 13976
rect 18354 13914 18388 13948
rect 13342 13822 13376 13856
rect 13342 13754 13376 13788
rect 13342 13686 13376 13720
rect 13342 13618 13376 13652
rect 13342 13550 13376 13584
rect 13342 13482 13376 13516
rect 18354 13846 18388 13880
rect 18354 13778 18388 13812
rect 18354 13710 18388 13744
rect 18354 13642 18388 13676
rect 18354 13574 18388 13608
rect 18354 13506 18388 13540
rect 13342 13414 13376 13448
rect 13342 13346 13376 13380
rect 13462 13346 13496 13458
rect 14018 13346 14052 13460
rect 15130 13346 15164 13439
rect 18354 13438 18388 13472
rect 15792 13346 15826 13420
rect 16452 13346 16486 13420
rect 17670 13346 17704 13420
rect 18226 13346 18260 13420
rect 18354 13370 18388 13404
rect 13376 13312 13522 13346
rect 13342 13292 13522 13312
rect 13897 13292 14059 13346
rect 14530 13292 14692 13346
rect 15125 13292 15287 13346
rect 15785 13292 15947 13346
rect 16335 13292 16497 13346
rect 17004 13292 17166 13346
rect 17619 13292 17781 13346
rect 18210 13336 18354 13346
rect 18210 13302 18388 13336
rect 18210 13292 18354 13302
rect 13342 13278 13376 13292
rect 13342 13210 13376 13244
rect 18354 13234 18388 13268
rect 14680 13210 16668 13212
rect 13288 13176 13366 13210
rect 13400 13176 13434 13210
rect 13468 13176 13502 13210
rect 13536 13176 13570 13210
rect 13604 13176 13638 13210
rect 13672 13176 13706 13210
rect 13740 13176 13774 13210
rect 13808 13176 13842 13210
rect 13876 13176 13910 13210
rect 13944 13176 13978 13210
rect 14012 13176 14046 13210
rect 14080 13176 14114 13210
rect 14148 13176 14182 13210
rect 14216 13176 14250 13210
rect 14284 13176 14318 13210
rect 14352 13176 14386 13210
rect 14420 13176 14454 13210
rect 14488 13176 14522 13210
rect 14556 13176 14590 13210
rect 14624 13176 14658 13210
rect 14692 13176 14726 13210
rect 14760 13176 14794 13210
rect 14828 13176 14862 13210
rect 14896 13176 14930 13210
rect 14964 13176 14998 13210
rect 15032 13176 15066 13210
rect 15100 13176 15134 13210
rect 15168 13176 15202 13210
rect 15236 13176 15270 13210
rect 15304 13176 15338 13210
rect 15372 13176 15406 13210
rect 15440 13176 15474 13210
rect 15508 13176 15542 13210
rect 15576 13176 15610 13210
rect 15644 13176 15678 13210
rect 15712 13176 15746 13210
rect 15780 13176 15889 13210
rect 15923 13176 15957 13210
rect 15991 13176 16025 13210
rect 16059 13176 16093 13210
rect 16127 13176 16161 13210
rect 16195 13176 16229 13210
rect 16263 13176 16297 13210
rect 16331 13176 16365 13210
rect 16399 13176 16433 13210
rect 16467 13176 16501 13210
rect 16535 13176 16569 13210
rect 16603 13176 16637 13210
rect 16671 13176 16705 13210
rect 16739 13176 16773 13210
rect 16807 13176 16841 13210
rect 16875 13176 16909 13210
rect 16943 13176 16977 13210
rect 17011 13176 17045 13210
rect 17079 13176 17113 13210
rect 17147 13176 17181 13210
rect 17215 13176 17249 13210
rect 17283 13176 17317 13210
rect 17351 13176 17385 13210
rect 17419 13176 17453 13210
rect 17487 13176 17521 13210
rect 17555 13176 17589 13210
rect 17623 13176 17657 13210
rect 17691 13176 17725 13210
rect 17759 13176 17793 13210
rect 17827 13176 17861 13210
rect 17895 13176 17929 13210
rect 17963 13176 17997 13210
rect 18031 13176 18065 13210
rect 18099 13176 18133 13210
rect 18167 13176 18201 13210
rect 18235 13176 18269 13210
rect 18303 13200 18354 13210
rect 18303 13176 18388 13200
rect 13254 13142 13288 13176
rect 13254 13074 13288 13108
rect 13254 13006 13288 13040
rect 13534 12975 13734 13176
rect 14680 12972 16668 13176
rect 13254 12938 13288 12972
rect 13254 12870 13288 12904
rect 13254 12802 13288 12836
rect 13254 12734 13288 12768
rect 13388 12814 13458 12830
rect 13667 12823 13895 12857
rect 13388 12780 13408 12814
rect 13442 12780 13458 12814
rect 13388 12762 13458 12780
rect 13254 12666 13288 12700
rect 13254 12598 13288 12632
rect 13254 12530 13288 12564
rect 13254 12462 13288 12496
rect 13254 12394 13288 12428
rect 13254 12326 13288 12360
rect 13254 12258 13288 12292
rect 13254 12190 13288 12224
rect 13254 12122 13288 12156
rect 13254 12054 13288 12088
rect 13254 11986 13288 12020
rect 13254 11918 13288 11952
rect 13254 11850 13288 11884
rect 13254 11782 13288 11816
rect 11446 11730 11480 11764
rect 11446 11662 11480 11696
rect 11446 11594 11480 11628
rect 11446 11526 11480 11560
rect 11446 11458 11480 11492
rect 11996 11762 12032 11778
rect 11996 11728 11997 11762
rect 12031 11728 12032 11762
rect 11996 11690 12032 11728
rect 11996 11656 11997 11690
rect 12031 11656 12032 11690
rect 11996 11618 12032 11656
rect 11996 11584 11997 11618
rect 12031 11584 12032 11618
rect 11996 11546 12032 11584
rect 11996 11512 11997 11546
rect 12031 11512 12032 11546
rect 11996 11474 12032 11512
rect 11996 11440 11997 11474
rect 12031 11440 12032 11474
rect 11996 11424 12032 11440
rect 13254 11714 13288 11748
rect 13254 11646 13288 11680
rect 13254 11578 13288 11612
rect 13254 11510 13288 11544
rect 13254 11442 13288 11476
rect 11446 11390 11480 11424
rect 11446 11322 11480 11356
rect 11446 11254 11480 11288
rect 13254 11374 13288 11408
rect 13254 11306 13288 11340
rect 13254 11238 13288 11272
rect 11480 11220 11635 11232
rect 11446 11186 11635 11220
rect 11480 11178 11635 11186
rect 11962 11178 13023 11232
rect 13089 11204 13254 11232
rect 13089 11178 13288 11204
rect 11446 11118 11480 11152
rect 13254 11170 13288 11178
rect 13254 11094 13288 11136
rect 11480 11084 11530 11094
rect 11446 11060 11530 11084
rect 11564 11060 11598 11094
rect 11632 11060 11666 11094
rect 11700 11060 11734 11094
rect 11768 11060 11802 11094
rect 11836 11060 11870 11094
rect 11904 11060 11938 11094
rect 11972 11060 12006 11094
rect 12040 11060 12074 11094
rect 12108 11060 12142 11094
rect 12176 11060 12210 11094
rect 12244 11060 12278 11094
rect 12312 11060 12346 11094
rect 12380 11060 12414 11094
rect 12448 11060 12482 11094
rect 12516 11060 12550 11094
rect 12584 11060 12618 11094
rect 12652 11060 12686 11094
rect 12720 11060 12754 11094
rect 12788 11060 12822 11094
rect 12856 11060 12890 11094
rect 12924 11060 12958 11094
rect 12992 11060 13026 11094
rect 13060 11060 13094 11094
rect 13128 11060 13162 11094
rect 13196 11060 13230 11094
rect 13264 11060 13288 11094
rect 11446 10104 11652 11060
rect 14248 10498 14870 10930
rect 10248 7400 10318 9140
rect 10646 7390 10716 9212
rect 11536 7384 11606 9206
rect 11934 7390 12004 9212
rect 12826 7390 12896 9212
rect 14248 9058 14530 10072
rect 14248 8200 14870 8632
rect 12974 6772 13780 7204
rect 15338 6436 15620 7204
rect 12936 6336 15620 6436
<< viali >>
rect 9617 37466 9633 37500
rect 9633 37466 9651 37500
rect 9689 37466 9701 37500
rect 9701 37466 9723 37500
rect 9761 37466 9769 37500
rect 9769 37466 9795 37500
rect 9833 37466 9837 37500
rect 9837 37466 9867 37500
rect 9905 37466 9939 37500
rect 9977 37466 10007 37500
rect 10007 37466 10011 37500
rect 10049 37466 10075 37500
rect 10075 37466 10083 37500
rect 10121 37466 10143 37500
rect 10143 37466 10155 37500
rect 10193 37466 10211 37500
rect 10211 37466 10227 37500
rect 10358 37466 10374 37500
rect 10374 37466 10392 37500
rect 10430 37466 10442 37500
rect 10442 37466 10464 37500
rect 10502 37466 10510 37500
rect 10510 37466 10536 37500
rect 10574 37466 10578 37500
rect 10578 37466 10608 37500
rect 10646 37466 10680 37500
rect 10718 37466 10748 37500
rect 10748 37466 10752 37500
rect 10790 37466 10816 37500
rect 10816 37466 10824 37500
rect 10862 37466 10884 37500
rect 10884 37466 10896 37500
rect 10934 37466 10952 37500
rect 10952 37466 10968 37500
rect 11018 37466 11034 37500
rect 11034 37466 11052 37500
rect 11090 37466 11102 37500
rect 11102 37466 11124 37500
rect 11162 37466 11170 37500
rect 11170 37466 11196 37500
rect 11234 37466 11238 37500
rect 11238 37466 11268 37500
rect 11306 37466 11340 37500
rect 11378 37466 11408 37500
rect 11408 37466 11412 37500
rect 11450 37466 11476 37500
rect 11476 37466 11484 37500
rect 11522 37466 11544 37500
rect 11544 37466 11556 37500
rect 11594 37466 11612 37500
rect 11612 37466 11628 37500
rect 11674 37466 11690 37500
rect 11690 37466 11708 37500
rect 11746 37466 11758 37500
rect 11758 37466 11780 37500
rect 11818 37466 11826 37500
rect 11826 37466 11852 37500
rect 11890 37466 11894 37500
rect 11894 37466 11924 37500
rect 11962 37466 11996 37500
rect 12034 37466 12064 37500
rect 12064 37466 12068 37500
rect 12106 37466 12132 37500
rect 12132 37466 12140 37500
rect 12178 37466 12200 37500
rect 12200 37466 12212 37500
rect 12250 37466 12268 37500
rect 12268 37466 12284 37500
rect 12347 37466 12363 37500
rect 12363 37466 12381 37500
rect 12419 37466 12431 37500
rect 12431 37466 12453 37500
rect 12491 37466 12499 37500
rect 12499 37466 12525 37500
rect 12563 37466 12567 37500
rect 12567 37466 12597 37500
rect 12635 37466 12669 37500
rect 12707 37466 12737 37500
rect 12737 37466 12741 37500
rect 12779 37466 12805 37500
rect 12805 37466 12813 37500
rect 12851 37466 12873 37500
rect 12873 37466 12885 37500
rect 12923 37466 12941 37500
rect 12941 37466 12957 37500
rect 13020 37466 13036 37500
rect 13036 37466 13054 37500
rect 13092 37466 13104 37500
rect 13104 37466 13126 37500
rect 13164 37466 13172 37500
rect 13172 37466 13198 37500
rect 13236 37466 13240 37500
rect 13240 37466 13270 37500
rect 13308 37466 13342 37500
rect 13380 37466 13410 37500
rect 13410 37466 13414 37500
rect 13452 37466 13478 37500
rect 13478 37466 13486 37500
rect 13524 37466 13546 37500
rect 13546 37466 13558 37500
rect 13596 37466 13614 37500
rect 13614 37466 13630 37500
rect 13680 37466 13696 37500
rect 13696 37466 13714 37500
rect 13752 37466 13764 37500
rect 13764 37466 13786 37500
rect 13824 37466 13832 37500
rect 13832 37466 13858 37500
rect 13896 37466 13900 37500
rect 13900 37466 13930 37500
rect 13968 37466 14002 37500
rect 14040 37466 14070 37500
rect 14070 37466 14074 37500
rect 14112 37466 14138 37500
rect 14138 37466 14146 37500
rect 14184 37466 14206 37500
rect 14206 37466 14218 37500
rect 14256 37466 14274 37500
rect 14274 37466 14290 37500
rect 19127 37448 19143 37482
rect 19143 37448 19161 37482
rect 19199 37448 19211 37482
rect 19211 37448 19233 37482
rect 19271 37448 19279 37482
rect 19279 37448 19305 37482
rect 19343 37448 19347 37482
rect 19347 37448 19377 37482
rect 19415 37448 19449 37482
rect 19487 37448 19517 37482
rect 19517 37448 19521 37482
rect 19559 37448 19585 37482
rect 19585 37448 19593 37482
rect 19631 37448 19653 37482
rect 19653 37448 19665 37482
rect 19703 37448 19721 37482
rect 19721 37448 19737 37482
rect 19800 37448 19816 37482
rect 19816 37448 19834 37482
rect 19872 37448 19884 37482
rect 19884 37448 19906 37482
rect 19944 37448 19952 37482
rect 19952 37448 19978 37482
rect 20016 37448 20020 37482
rect 20020 37448 20050 37482
rect 20088 37448 20122 37482
rect 20160 37448 20190 37482
rect 20190 37448 20194 37482
rect 20232 37448 20258 37482
rect 20258 37448 20266 37482
rect 20304 37448 20326 37482
rect 20326 37448 20338 37482
rect 20376 37448 20394 37482
rect 20394 37448 20410 37482
rect 20475 37448 20489 37482
rect 20489 37448 20509 37482
rect 20547 37448 20557 37482
rect 20557 37448 20581 37482
rect 20619 37448 20625 37482
rect 20625 37448 20653 37482
rect 20691 37448 20693 37482
rect 20693 37448 20725 37482
rect 20763 37448 20795 37482
rect 20795 37448 20797 37482
rect 20835 37448 20863 37482
rect 20863 37448 20869 37482
rect 20907 37448 20931 37482
rect 20931 37448 20941 37482
rect 20979 37448 20999 37482
rect 20999 37448 21013 37482
rect 21078 37448 21094 37482
rect 21094 37448 21112 37482
rect 21150 37448 21162 37482
rect 21162 37448 21184 37482
rect 21222 37448 21230 37482
rect 21230 37448 21256 37482
rect 21294 37448 21298 37482
rect 21298 37448 21328 37482
rect 21366 37448 21400 37482
rect 21438 37448 21468 37482
rect 21468 37448 21472 37482
rect 21510 37448 21536 37482
rect 21536 37448 21544 37482
rect 21582 37448 21604 37482
rect 21604 37448 21616 37482
rect 21654 37448 21672 37482
rect 21672 37448 21688 37482
rect 21751 37448 21767 37482
rect 21767 37448 21785 37482
rect 21823 37448 21835 37482
rect 21835 37448 21857 37482
rect 21895 37448 21903 37482
rect 21903 37448 21929 37482
rect 21967 37448 21971 37482
rect 21971 37448 22001 37482
rect 22039 37448 22073 37482
rect 22111 37448 22141 37482
rect 22141 37448 22145 37482
rect 22183 37448 22209 37482
rect 22209 37448 22217 37482
rect 22255 37448 22277 37482
rect 22277 37448 22289 37482
rect 22327 37448 22345 37482
rect 22345 37448 22361 37482
rect 22424 37448 22440 37482
rect 22440 37448 22458 37482
rect 22496 37448 22508 37482
rect 22508 37448 22530 37482
rect 22568 37448 22576 37482
rect 22576 37448 22602 37482
rect 22640 37448 22644 37482
rect 22644 37448 22674 37482
rect 22712 37448 22746 37482
rect 22784 37448 22814 37482
rect 22814 37448 22818 37482
rect 22856 37448 22882 37482
rect 22882 37448 22890 37482
rect 22928 37448 22950 37482
rect 22950 37448 22962 37482
rect 23000 37448 23018 37482
rect 23018 37448 23034 37482
rect 9638 34532 9672 34566
rect 9714 34532 9748 34566
rect 9790 34532 9824 34566
rect 9866 34532 9900 34566
rect 9942 34532 9976 34566
rect 10018 34532 10052 34566
rect 10095 34532 10129 34566
rect 10172 34532 10206 34566
rect 10400 34532 10434 34566
rect 10476 34532 10510 34566
rect 10552 34532 10586 34566
rect 10628 34532 10662 34566
rect 10704 34532 10738 34566
rect 10780 34532 10814 34566
rect 10857 34532 10891 34566
rect 10934 34532 10968 34566
rect 11056 34532 11090 34566
rect 11132 34532 11166 34566
rect 11208 34532 11242 34566
rect 11284 34532 11318 34566
rect 11360 34532 11394 34566
rect 11436 34532 11470 34566
rect 11513 34532 11547 34566
rect 11590 34532 11624 34566
rect 11712 34532 11746 34566
rect 11789 34532 11823 34566
rect 11866 34532 11900 34566
rect 11942 34532 11976 34566
rect 12018 34532 12052 34566
rect 12094 34532 12128 34566
rect 12170 34532 12204 34566
rect 12246 34532 12280 34566
rect 12368 34532 12402 34566
rect 12444 34532 12478 34566
rect 12520 34532 12554 34566
rect 12596 34532 12630 34566
rect 12672 34532 12706 34566
rect 12748 34532 12782 34566
rect 12825 34532 12859 34566
rect 12902 34532 12936 34566
rect 13024 34532 13058 34566
rect 13101 34532 13135 34566
rect 13178 34532 13212 34566
rect 13254 34532 13288 34566
rect 13330 34532 13364 34566
rect 13406 34532 13440 34566
rect 13482 34532 13516 34566
rect 13558 34532 13592 34566
rect 13680 34532 13714 34566
rect 13757 34532 13791 34566
rect 13834 34532 13868 34566
rect 13910 34532 13944 34566
rect 13986 34532 14020 34566
rect 14062 34532 14096 34566
rect 14138 34532 14172 34566
rect 14214 34532 14248 34566
rect 9289 34364 9323 34398
rect 9836 34147 9870 34181
rect 9970 34147 10004 34181
rect 10092 34147 10126 34181
rect 10226 34147 10260 34181
rect 9667 34054 9701 34068
rect 9667 34034 9701 34054
rect 9667 33986 9701 33996
rect 8606 33610 8640 33644
rect 9667 33962 9701 33986
rect 9667 33918 9701 33924
rect 9667 33890 9701 33918
rect 9667 33850 9701 33852
rect 9667 33818 9701 33850
rect 9667 33748 9701 33780
rect 9667 33746 9701 33748
rect 9667 33680 9701 33708
rect 9667 33674 9701 33680
rect 9667 33612 9701 33636
rect 9667 33602 9701 33612
rect 9667 33544 9701 33564
rect 9667 33530 9701 33544
rect 8045 33354 8079 33388
rect 10966 34147 11000 34181
rect 11100 34147 11134 34181
rect 11222 34147 11256 34181
rect 11356 34147 11390 34181
rect 11525 34054 11559 34068
rect 11525 34034 11559 34054
rect 11525 33986 11559 33996
rect 11525 33962 11559 33986
rect 11525 33918 11559 33924
rect 11525 33890 11559 33918
rect 11525 33850 11559 33852
rect 11525 33818 11559 33850
rect 11525 33748 11559 33780
rect 11525 33746 11559 33748
rect 11525 33680 11559 33708
rect 11525 33674 11559 33680
rect 11525 33612 11559 33636
rect 11525 33602 11559 33612
rect 11525 33544 11559 33564
rect 11525 33530 11559 33544
rect 9836 33417 9870 33451
rect 9970 33417 10004 33451
rect 10092 33417 10126 33451
rect 10226 33417 10260 33451
rect 10348 33417 10382 33451
rect 10482 33417 10516 33451
rect 10710 33417 10744 33451
rect 10844 33417 10878 33451
rect 10966 33417 11000 33451
rect 11100 33417 11134 33451
rect 11222 33417 11256 33451
rect 11356 33417 11390 33451
rect 7521 33138 7555 33172
rect 11998 34204 12002 34238
rect 12002 34204 12032 34238
rect 12070 34204 12104 34238
rect 12142 34204 12172 34238
rect 12172 34204 12176 34238
rect 12258 34204 12262 34238
rect 12262 34204 12292 34238
rect 12330 34204 12364 34238
rect 12402 34204 12432 34238
rect 12432 34204 12436 34238
rect 12499 34204 12505 34238
rect 12505 34204 12533 34238
rect 12571 34204 12573 34238
rect 12573 34204 12605 34238
rect 12643 34204 12675 34238
rect 12675 34204 12677 34238
rect 12715 34204 12743 34238
rect 12743 34204 12749 34238
rect 13137 34186 13153 34220
rect 13153 34186 13171 34220
rect 13209 34186 13221 34220
rect 13221 34186 13243 34220
rect 13281 34186 13289 34220
rect 13289 34186 13315 34220
rect 13353 34186 13357 34220
rect 13357 34186 13387 34220
rect 13425 34186 13459 34220
rect 13497 34186 13527 34220
rect 13527 34186 13531 34220
rect 13569 34186 13595 34220
rect 13595 34186 13603 34220
rect 13641 34186 13663 34220
rect 13663 34186 13675 34220
rect 13713 34186 13731 34220
rect 13731 34186 13747 34220
rect 13911 34186 13927 34220
rect 13927 34186 13945 34220
rect 13983 34186 13995 34220
rect 13995 34186 14017 34220
rect 14055 34186 14063 34220
rect 14063 34186 14089 34220
rect 14127 34186 14131 34220
rect 14131 34186 14161 34220
rect 14199 34186 14233 34220
rect 14271 34186 14301 34220
rect 14301 34186 14305 34220
rect 14343 34186 14369 34220
rect 14369 34186 14377 34220
rect 14415 34186 14437 34220
rect 14437 34186 14449 34220
rect 14487 34186 14505 34220
rect 14505 34186 14521 34220
rect 12024 33332 12058 33366
rect 12158 33332 12192 33366
rect 12280 33332 12314 33366
rect 12414 33332 12448 33366
rect 12536 33332 12570 33366
rect 12670 33332 12704 33366
rect 19348 33848 19382 33882
rect 13158 33349 13192 33383
rect 13234 33349 13268 33383
rect 13310 33349 13344 33383
rect 13386 33349 13420 33383
rect 13462 33349 13496 33383
rect 13538 33349 13572 33383
rect 13615 33349 13649 33383
rect 13692 33349 13726 33383
rect 13936 33349 13970 33383
rect 14012 33349 14046 33383
rect 14088 33349 14122 33383
rect 14164 33349 14198 33383
rect 14240 33349 14274 33383
rect 14316 33349 14350 33383
rect 14393 33349 14427 33383
rect 14470 33349 14504 33383
rect 21855 33392 22249 33642
rect 23374 33392 23768 33642
rect 9096 33136 9130 33170
rect 21855 33062 22249 33312
rect 23374 33062 23768 33312
rect 7389 32959 7423 32993
rect 8542 32912 8576 32946
rect 9642 32876 9650 32910
rect 9650 32876 9676 32910
rect 9714 32876 9718 32910
rect 9718 32876 9748 32910
rect 9786 32876 9820 32910
rect 9858 32876 9888 32910
rect 9888 32876 9892 32910
rect 9930 32876 9956 32910
rect 9956 32876 9964 32910
rect 10038 32876 10044 32910
rect 10044 32876 10072 32910
rect 10110 32876 10112 32910
rect 10112 32876 10144 32910
rect 10182 32876 10214 32910
rect 10214 32876 10216 32910
rect 10254 32876 10282 32910
rect 10282 32876 10288 32910
rect 10394 32876 10400 32910
rect 10400 32876 10428 32910
rect 10466 32876 10468 32910
rect 10468 32876 10500 32910
rect 10538 32876 10570 32910
rect 10570 32876 10572 32910
rect 10610 32876 10638 32910
rect 10638 32876 10644 32910
rect 10735 32876 10743 32910
rect 10743 32876 10769 32910
rect 10807 32876 10811 32910
rect 10811 32876 10841 32910
rect 10879 32876 10913 32910
rect 10951 32876 10981 32910
rect 10981 32876 10985 32910
rect 11023 32876 11049 32910
rect 11049 32876 11057 32910
rect 11511 32896 11545 32930
rect 11584 32896 11618 32930
rect 11657 32896 11691 32930
rect 11729 32896 11763 32930
rect 11801 32896 11835 32930
rect 11873 32896 11907 32930
rect 11945 32896 11979 32930
rect 12067 32896 12101 32930
rect 12140 32896 12174 32930
rect 12213 32896 12247 32930
rect 12285 32896 12319 32930
rect 12357 32896 12391 32930
rect 12429 32896 12463 32930
rect 12501 32896 12535 32930
rect 12623 32896 12657 32930
rect 12695 32896 12729 32930
rect 12767 32896 12801 32930
rect 12839 32896 12873 32930
rect 12911 32896 12945 32930
rect 12984 32896 13018 32930
rect 13057 32896 13091 32930
rect 13285 32896 13319 32930
rect 13357 32896 13391 32930
rect 13429 32896 13463 32930
rect 13501 32896 13535 32930
rect 13573 32896 13607 32930
rect 13646 32896 13680 32930
rect 13719 32896 13753 32930
rect 13841 32896 13875 32930
rect 13914 32896 13948 32930
rect 13987 32896 14021 32930
rect 14059 32896 14093 32930
rect 14131 32896 14165 32930
rect 14203 32896 14237 32930
rect 14275 32896 14309 32930
rect 8886 32676 8920 32710
rect 11091 32544 11125 32578
rect 21855 32732 22249 32982
rect 23374 32732 23768 32982
rect 21855 32400 22249 32650
rect 23374 32400 23768 32650
rect 21855 32072 22249 32322
rect 23374 32072 23768 32322
rect 11491 31678 11503 31712
rect 11503 31678 11525 31712
rect 11563 31678 11571 31712
rect 11571 31678 11597 31712
rect 11635 31678 11639 31712
rect 11639 31678 11669 31712
rect 11707 31678 11741 31712
rect 11779 31678 11809 31712
rect 11809 31678 11813 31712
rect 11851 31678 11877 31712
rect 11877 31678 11885 31712
rect 11923 31678 11945 31712
rect 11945 31678 11957 31712
rect 12051 31678 12063 31712
rect 12063 31678 12085 31712
rect 12123 31678 12131 31712
rect 12131 31678 12157 31712
rect 12195 31678 12199 31712
rect 12199 31678 12229 31712
rect 12267 31678 12301 31712
rect 12339 31678 12369 31712
rect 12369 31678 12373 31712
rect 12411 31678 12437 31712
rect 12437 31678 12445 31712
rect 12483 31678 12505 31712
rect 12505 31678 12517 31712
rect 12592 31678 12606 31712
rect 12606 31678 12626 31712
rect 12664 31678 12674 31712
rect 12674 31678 12698 31712
rect 12736 31678 12742 31712
rect 12742 31678 12770 31712
rect 12808 31678 12810 31712
rect 12810 31678 12842 31712
rect 12880 31678 12912 31712
rect 12912 31678 12914 31712
rect 12952 31678 12980 31712
rect 12980 31678 12986 31712
rect 13024 31678 13048 31712
rect 13048 31678 13058 31712
rect 13096 31678 13116 31712
rect 13116 31678 13130 31712
rect 13246 31678 13260 31712
rect 13260 31678 13280 31712
rect 13318 31678 13328 31712
rect 13328 31678 13352 31712
rect 13390 31678 13396 31712
rect 13396 31678 13424 31712
rect 13462 31678 13464 31712
rect 13464 31678 13496 31712
rect 13534 31678 13566 31712
rect 13566 31678 13568 31712
rect 13606 31678 13634 31712
rect 13634 31678 13640 31712
rect 13678 31678 13702 31712
rect 13702 31678 13712 31712
rect 13750 31678 13770 31712
rect 13770 31678 13784 31712
rect 13863 31678 13875 31712
rect 13875 31678 13897 31712
rect 13935 31678 13943 31712
rect 13943 31678 13969 31712
rect 14007 31678 14011 31712
rect 14011 31678 14041 31712
rect 14079 31678 14113 31712
rect 14151 31678 14181 31712
rect 14181 31678 14185 31712
rect 14223 31678 14249 31712
rect 14249 31678 14257 31712
rect 14295 31678 14317 31712
rect 14317 31678 14329 31712
rect 21855 31742 22249 31992
rect 23374 31742 23768 31992
rect 9690 31312 9724 31346
rect 9768 31312 9802 31346
rect 9846 31312 9880 31346
rect 9924 31312 9958 31346
rect 10046 31312 10080 31346
rect 10124 31312 10158 31346
rect 10202 31312 10236 31346
rect 10280 31312 10314 31346
rect 10402 31312 10436 31346
rect 10480 31312 10514 31346
rect 10558 31312 10592 31346
rect 10636 31312 10670 31346
rect 10758 31312 10792 31346
rect 10836 31312 10870 31346
rect 10914 31312 10948 31346
rect 10992 31312 11026 31346
rect 21855 31412 22249 31662
rect 23374 31412 23768 31662
rect 9690 31128 9724 31162
rect 9768 31128 9802 31162
rect 9846 31128 9880 31162
rect 9924 31128 9958 31162
rect 10046 31128 10080 31162
rect 10124 31128 10158 31162
rect 10202 31128 10236 31162
rect 10280 31128 10314 31162
rect 10402 31128 10436 31162
rect 10480 31128 10514 31162
rect 10558 31128 10592 31162
rect 10636 31128 10670 31162
rect 10758 31128 10792 31162
rect 10836 31128 10870 31162
rect 10914 31128 10948 31162
rect 10992 31128 11026 31162
rect 11396 31156 11430 31190
rect 12817 31198 12851 31232
rect 12889 31198 12923 31232
rect 12961 31198 12995 31232
rect 13033 31198 13067 31232
rect 13105 31198 13139 31232
rect 13177 31198 13211 31232
rect 14076 31198 14110 31232
rect 14148 31198 14182 31232
rect 14220 31198 14254 31232
rect 14292 31198 14326 31232
rect 14364 31198 14398 31232
rect 14436 31198 14470 31232
rect 9985 30125 10019 30138
rect 9985 30104 10019 30125
rect 9985 30057 10019 30066
rect 9985 30032 10019 30057
rect 9985 29989 10019 29994
rect 9985 29960 10019 29989
rect 9985 29921 10019 29922
rect 9985 29888 10019 29921
rect 9985 29819 10019 29850
rect 9985 29816 10019 29819
rect 21855 31082 22249 31332
rect 23374 31082 23768 31332
rect 9659 29564 9667 29598
rect 9667 29564 9693 29598
rect 9731 29564 9735 29598
rect 9735 29564 9765 29598
rect 9803 29564 9837 29598
rect 9875 29564 9905 29598
rect 9905 29564 9909 29598
rect 9947 29564 9973 29598
rect 9973 29564 9981 29598
rect 10072 29564 10078 29598
rect 10078 29564 10106 29598
rect 10144 29564 10146 29598
rect 10146 29564 10178 29598
rect 10216 29564 10248 29598
rect 10248 29564 10250 29598
rect 10288 29564 10316 29598
rect 10316 29564 10322 29598
rect 10411 29564 10417 29598
rect 10417 29564 10445 29598
rect 10483 29564 10485 29598
rect 10485 29564 10517 29598
rect 10555 29564 10587 29598
rect 10587 29564 10589 29598
rect 10627 29564 10655 29598
rect 10655 29564 10661 29598
rect 10735 29564 10743 29598
rect 10743 29564 10769 29598
rect 10807 29564 10811 29598
rect 10811 29564 10841 29598
rect 10879 29564 10913 29598
rect 10951 29564 10981 29598
rect 10981 29564 10985 29598
rect 11023 29564 11049 29598
rect 11049 29564 11057 29598
rect 10618 15234 10652 15268
rect 10057 14978 10091 15012
rect 9533 14762 9567 14796
rect 21360 15472 21394 15506
rect 11108 14760 11142 14794
rect 9401 14583 9435 14617
rect 10554 14536 10588 14570
rect 10898 14300 10932 14334
rect 13103 14168 13137 14202
rect 9191 12369 9297 12475
rect 13408 12780 13442 12814
rect 11997 11728 12031 11762
rect 11997 11656 12031 11690
rect 11997 11584 12031 11618
rect 11997 11512 12031 11546
rect 11997 11440 12031 11474
<< metal1 >>
rect 9571 37500 15288 37510
rect 9571 37466 9617 37500
rect 9651 37466 9689 37500
rect 9723 37466 9761 37500
rect 9795 37466 9833 37500
rect 9867 37466 9905 37500
rect 9939 37466 9977 37500
rect 10011 37466 10049 37500
rect 10083 37466 10121 37500
rect 10155 37466 10193 37500
rect 10227 37466 10358 37500
rect 10392 37466 10430 37500
rect 10464 37466 10502 37500
rect 10536 37466 10574 37500
rect 10608 37466 10646 37500
rect 10680 37466 10718 37500
rect 10752 37466 10790 37500
rect 10824 37466 10862 37500
rect 10896 37466 10934 37500
rect 10968 37466 11018 37500
rect 11052 37466 11090 37500
rect 11124 37466 11162 37500
rect 11196 37466 11234 37500
rect 11268 37466 11306 37500
rect 11340 37466 11378 37500
rect 11412 37466 11450 37500
rect 11484 37466 11522 37500
rect 11556 37466 11594 37500
rect 11628 37466 11674 37500
rect 11708 37466 11746 37500
rect 11780 37466 11818 37500
rect 11852 37466 11890 37500
rect 11924 37466 11962 37500
rect 11996 37466 12034 37500
rect 12068 37466 12106 37500
rect 12140 37466 12178 37500
rect 12212 37466 12250 37500
rect 12284 37466 12347 37500
rect 12381 37466 12419 37500
rect 12453 37466 12491 37500
rect 12525 37466 12563 37500
rect 12597 37466 12635 37500
rect 12669 37466 12707 37500
rect 12741 37466 12779 37500
rect 12813 37466 12851 37500
rect 12885 37466 12923 37500
rect 12957 37466 13020 37500
rect 13054 37466 13092 37500
rect 13126 37466 13164 37500
rect 13198 37466 13236 37500
rect 13270 37466 13308 37500
rect 13342 37466 13380 37500
rect 13414 37466 13452 37500
rect 13486 37466 13524 37500
rect 13558 37466 13596 37500
rect 13630 37466 13680 37500
rect 13714 37466 13752 37500
rect 13786 37466 13824 37500
rect 13858 37466 13896 37500
rect 13930 37466 13968 37500
rect 14002 37466 14040 37500
rect 14074 37466 14112 37500
rect 14146 37466 14184 37500
rect 14218 37466 14256 37500
rect 14290 37492 15288 37500
rect 14290 37482 23719 37492
rect 14290 37466 19127 37482
rect 9571 37456 19127 37466
rect 15234 37448 19127 37456
rect 19161 37448 19199 37482
rect 19233 37448 19271 37482
rect 19305 37448 19343 37482
rect 19377 37448 19415 37482
rect 19449 37448 19487 37482
rect 19521 37448 19559 37482
rect 19593 37448 19631 37482
rect 19665 37448 19703 37482
rect 19737 37448 19800 37482
rect 19834 37448 19872 37482
rect 19906 37448 19944 37482
rect 19978 37448 20016 37482
rect 20050 37448 20088 37482
rect 20122 37448 20160 37482
rect 20194 37448 20232 37482
rect 20266 37448 20304 37482
rect 20338 37448 20376 37482
rect 20410 37448 20475 37482
rect 20509 37448 20547 37482
rect 20581 37448 20619 37482
rect 20653 37448 20691 37482
rect 20725 37448 20763 37482
rect 20797 37448 20835 37482
rect 20869 37448 20907 37482
rect 20941 37448 20979 37482
rect 21013 37448 21078 37482
rect 21112 37448 21150 37482
rect 21184 37448 21222 37482
rect 21256 37448 21294 37482
rect 21328 37448 21366 37482
rect 21400 37448 21438 37482
rect 21472 37448 21510 37482
rect 21544 37448 21582 37482
rect 21616 37448 21654 37482
rect 21688 37448 21751 37482
rect 21785 37448 21823 37482
rect 21857 37448 21895 37482
rect 21929 37448 21967 37482
rect 22001 37448 22039 37482
rect 22073 37448 22111 37482
rect 22145 37448 22183 37482
rect 22217 37448 22255 37482
rect 22289 37448 22327 37482
rect 22361 37448 22424 37482
rect 22458 37448 22496 37482
rect 22530 37448 22568 37482
rect 22602 37448 22640 37482
rect 22674 37448 22712 37482
rect 22746 37448 22784 37482
rect 22818 37448 22856 37482
rect 22890 37448 22928 37482
rect 22962 37448 23000 37482
rect 23034 37448 23719 37482
rect 15234 37438 23719 37448
rect 18425 37436 18479 37438
rect 10990 36374 13654 36576
rect 5606 35987 5676 36020
rect 5606 35935 5614 35987
rect 5666 35935 5676 35987
rect 5606 35906 5676 35935
rect 5722 35758 5892 36180
rect 5944 35756 6114 36178
rect 6170 35756 6340 36178
rect 6394 35756 6564 36178
rect 6664 35900 7242 36020
rect 7576 35978 7676 36020
rect 7576 35926 7602 35978
rect 7654 35926 7676 35978
rect 7576 35906 7676 35926
rect 7142 35828 7242 35900
rect 7142 35776 7166 35828
rect 7218 35776 7242 35828
rect 7142 35766 7242 35776
rect 7600 34382 7654 35906
rect 10250 35898 14398 36100
rect 16090 35973 17402 36007
rect 19075 35962 20416 36020
rect 9622 34566 10984 34576
rect 9622 34532 9638 34566
rect 9672 34532 9714 34566
rect 9748 34532 9790 34566
rect 9824 34532 9866 34566
rect 9900 34532 9942 34566
rect 9976 34532 10018 34566
rect 10052 34532 10095 34566
rect 10129 34532 10172 34566
rect 10206 34532 10400 34566
rect 10434 34532 10476 34566
rect 10510 34532 10552 34566
rect 10586 34532 10628 34566
rect 10662 34532 10704 34566
rect 10738 34532 10780 34566
rect 10814 34532 10857 34566
rect 10891 34532 10934 34566
rect 10968 34532 10984 34566
rect 9622 34522 10984 34532
rect 11040 34566 13608 34576
rect 11040 34532 11056 34566
rect 11090 34532 11132 34566
rect 11166 34532 11208 34566
rect 11242 34532 11284 34566
rect 11318 34532 11360 34566
rect 11394 34532 11436 34566
rect 11470 34532 11513 34566
rect 11547 34532 11590 34566
rect 11624 34532 11712 34566
rect 11746 34532 11789 34566
rect 11823 34532 11866 34566
rect 11900 34532 11942 34566
rect 11976 34532 12018 34566
rect 12052 34532 12094 34566
rect 12128 34532 12170 34566
rect 12204 34532 12246 34566
rect 12280 34532 12368 34566
rect 12402 34532 12444 34566
rect 12478 34532 12520 34566
rect 12554 34532 12596 34566
rect 12630 34532 12672 34566
rect 12706 34532 12748 34566
rect 12782 34532 12825 34566
rect 12859 34532 12902 34566
rect 12936 34532 13024 34566
rect 13058 34532 13101 34566
rect 13135 34532 13178 34566
rect 13212 34532 13254 34566
rect 13288 34532 13330 34566
rect 13364 34532 13406 34566
rect 13440 34532 13482 34566
rect 13516 34532 13558 34566
rect 13592 34532 13608 34566
rect 11040 34522 13608 34532
rect 13664 34566 14600 34576
rect 13664 34532 13680 34566
rect 13714 34532 13757 34566
rect 13791 34532 13834 34566
rect 13868 34532 13910 34566
rect 13944 34532 13986 34566
rect 14020 34532 14062 34566
rect 14096 34532 14138 34566
rect 14172 34532 14214 34566
rect 14248 34532 14600 34566
rect 13664 34522 14600 34532
rect 15026 34522 15516 34576
rect 16391 34522 17123 34576
rect 9014 34409 9352 34448
rect 9014 34357 9029 34409
rect 9081 34398 9352 34409
rect 9081 34364 9289 34398
rect 9323 34364 9352 34398
rect 12356 34387 12558 34522
rect 16721 34441 16775 34522
rect 17490 34374 17570 34576
rect 17579 34532 17624 34576
rect 17749 34532 18613 34576
rect 17752 34522 18613 34532
rect 19302 34522 20088 34576
rect 20631 34522 20744 34576
rect 19734 34441 19788 34522
rect 9081 34357 9352 34364
rect 9014 34318 9352 34357
rect 16500 34334 17570 34374
rect 16500 34262 16762 34334
rect 11957 34238 12771 34248
rect 11957 34204 11998 34238
rect 12032 34204 12070 34238
rect 12104 34204 12142 34238
rect 12176 34204 12258 34238
rect 12292 34204 12330 34238
rect 12364 34204 12402 34238
rect 12436 34204 12499 34238
rect 12533 34204 12571 34238
rect 12605 34204 12643 34238
rect 12677 34204 12715 34238
rect 12749 34204 12771 34238
rect 11957 34194 12771 34204
rect 13091 34220 15868 34230
rect 9657 34181 11569 34191
rect 9657 34147 9836 34181
rect 9870 34147 9970 34181
rect 10004 34147 10092 34181
rect 10126 34147 10226 34181
rect 10260 34147 10966 34181
rect 11000 34147 11100 34181
rect 11134 34147 11222 34181
rect 11256 34147 11356 34181
rect 11390 34147 11569 34181
rect 13091 34186 13137 34220
rect 13171 34186 13209 34220
rect 13243 34186 13281 34220
rect 13315 34186 13353 34220
rect 13387 34186 13425 34220
rect 13459 34186 13497 34220
rect 13531 34186 13569 34220
rect 13603 34186 13641 34220
rect 13675 34186 13713 34220
rect 13747 34186 13911 34220
rect 13945 34186 13983 34220
rect 14017 34186 14055 34220
rect 14089 34186 14127 34220
rect 14161 34186 14199 34220
rect 14233 34186 14271 34220
rect 14305 34186 14343 34220
rect 14377 34186 14415 34220
rect 14449 34186 14487 34220
rect 14521 34186 15868 34220
rect 13091 34176 15868 34186
rect 9657 34137 11569 34147
rect 9657 34068 9711 34137
rect 9657 34034 9667 34068
rect 9701 34034 9711 34068
rect 9657 33996 9711 34034
rect 9657 33962 9667 33996
rect 9701 33962 9711 33996
rect 9657 33924 9711 33962
rect 9657 33890 9667 33924
rect 9701 33890 9711 33924
rect 9657 33852 9711 33890
rect 9657 33818 9667 33852
rect 9701 33818 9711 33852
rect 9657 33780 9711 33818
rect 9657 33746 9667 33780
rect 9701 33746 9711 33780
rect 9657 33708 9711 33746
rect 9657 33674 9667 33708
rect 9701 33674 9711 33708
rect 8583 33654 8659 33663
rect 8583 33602 8596 33654
rect 8648 33602 8659 33654
rect 8583 33591 8659 33602
rect 9657 33636 9711 33674
rect 9657 33602 9667 33636
rect 9701 33602 9711 33636
rect 9657 33564 9711 33602
rect 8864 33547 8928 33552
rect 7909 33545 9021 33547
rect 7909 33493 8870 33545
rect 8922 33493 9021 33545
rect 9657 33530 9667 33564
rect 9701 33530 9711 33564
rect 8864 33488 8928 33493
rect 9657 33461 9711 33530
rect 11515 34068 11569 34137
rect 11515 34034 11525 34068
rect 11559 34034 11569 34068
rect 11515 33996 11569 34034
rect 11515 33962 11525 33996
rect 11559 33962 11569 33996
rect 11515 33924 11569 33962
rect 11515 33890 11525 33924
rect 11559 33890 11569 33924
rect 12356 33903 12558 34036
rect 11515 33852 11569 33890
rect 11515 33818 11525 33852
rect 11559 33818 11569 33852
rect 11515 33780 11569 33818
rect 11515 33746 11525 33780
rect 11559 33746 11569 33780
rect 11515 33708 11569 33746
rect 11515 33674 11525 33708
rect 11559 33674 11569 33708
rect 12236 33701 12748 33903
rect 15028 33868 16742 33880
rect 15028 33708 16762 33868
rect 16814 33858 17420 34290
rect 17462 33858 18068 34290
rect 18110 33858 18716 34290
rect 18774 34261 19024 34272
rect 18774 33889 18777 34261
rect 19021 34194 19024 34261
rect 19021 33992 19244 34194
rect 21373 34193 21427 34576
rect 21665 34522 23368 34576
rect 19347 33993 21427 34193
rect 19021 33889 19024 33992
rect 18774 33878 19024 33889
rect 19336 33882 19394 33896
rect 19336 33848 19348 33882
rect 19382 33848 19394 33882
rect 11515 33636 11569 33674
rect 11515 33602 11525 33636
rect 11559 33602 11569 33636
rect 11515 33564 11569 33602
rect 11515 33530 11525 33564
rect 11559 33530 11569 33564
rect 11515 33461 11569 33530
rect 9657 33451 10276 33461
rect 9657 33417 9836 33451
rect 9870 33417 9970 33451
rect 10004 33417 10092 33451
rect 10126 33417 10226 33451
rect 10260 33417 10276 33451
rect 9657 33407 10276 33417
rect 10332 33451 10894 33461
rect 10332 33417 10348 33451
rect 10382 33417 10482 33451
rect 10516 33417 10710 33451
rect 10744 33417 10844 33451
rect 10878 33417 10894 33451
rect 10332 33407 10894 33417
rect 10950 33451 11569 33461
rect 10950 33417 10966 33451
rect 11000 33417 11100 33451
rect 11134 33417 11222 33451
rect 11256 33417 11356 33451
rect 11390 33417 11569 33451
rect 10950 33407 11569 33417
rect 7050 33180 7104 33396
rect 8034 33388 8094 33406
rect 15028 33393 15172 33708
rect 19336 33706 19394 33848
rect 7776 33354 8045 33388
rect 8079 33354 8094 33388
rect 13142 33383 13742 33393
rect 7776 33352 8094 33354
rect 7498 33188 7584 33198
rect 7498 33180 7590 33188
rect 7050 33128 7512 33180
rect 7564 33128 7590 33180
rect 7050 32622 7104 33128
rect 7498 33120 7590 33128
rect 7498 33116 7584 33120
rect 7692 33093 7802 33352
rect 8034 33340 8094 33352
rect 12008 33366 12720 33376
rect 12008 33332 12024 33366
rect 12058 33332 12158 33366
rect 12192 33332 12280 33366
rect 12314 33332 12414 33366
rect 12448 33332 12536 33366
rect 12570 33332 12670 33366
rect 12704 33332 12720 33366
rect 13142 33349 13158 33383
rect 13192 33349 13234 33383
rect 13268 33349 13310 33383
rect 13344 33349 13386 33383
rect 13420 33349 13462 33383
rect 13496 33349 13538 33383
rect 13572 33349 13615 33383
rect 13649 33349 13692 33383
rect 13726 33349 13742 33383
rect 13142 33339 13742 33349
rect 13920 33383 15176 33393
rect 13920 33349 13936 33383
rect 13970 33349 14012 33383
rect 14046 33349 14088 33383
rect 14122 33349 14164 33383
rect 14198 33349 14240 33383
rect 14274 33349 14316 33383
rect 14350 33349 14393 33383
rect 14427 33349 14470 33383
rect 14504 33349 15176 33383
rect 13920 33339 15176 33349
rect 12008 33322 12720 33332
rect 19552 33300 20138 33722
rect 20200 33300 20786 33722
rect 20848 33300 21434 33722
rect 21502 33687 21752 33698
rect 21502 33426 21505 33687
rect 21496 33315 21505 33426
rect 21749 33426 21752 33687
rect 21836 33642 22268 33658
rect 21749 33315 21758 33426
rect 21836 33392 21855 33642
rect 22249 33392 22268 33642
rect 21836 33312 22268 33392
rect 23361 33642 23782 33648
rect 23361 33392 23374 33642
rect 23768 33392 23782 33642
rect 23361 33386 23782 33392
rect 9256 33184 9356 33226
rect 9062 33180 9356 33184
rect 9062 33170 9288 33180
rect 9062 33136 9096 33170
rect 9130 33136 9288 33170
rect 9062 33128 9288 33136
rect 9340 33128 9356 33180
rect 9062 33120 9356 33128
rect 7366 33002 7446 33024
rect 7366 32950 7380 33002
rect 7432 32950 7446 33002
rect 7692 32991 7901 33093
rect 9256 33090 9356 33120
rect 7692 32987 7802 32991
rect 7692 32964 7726 32987
rect 7366 32934 7446 32950
rect 8528 32950 8592 32962
rect 8528 32898 8534 32950
rect 8586 32898 8592 32950
rect 11274 32930 11995 32940
rect 11274 32920 11511 32930
rect 8528 32892 8592 32898
rect 9623 32910 11511 32920
rect 9623 32876 9642 32910
rect 9676 32876 9714 32910
rect 9748 32876 9786 32910
rect 9820 32876 9858 32910
rect 9892 32876 9930 32910
rect 9964 32876 10038 32910
rect 10072 32876 10110 32910
rect 10144 32876 10182 32910
rect 10216 32876 10254 32910
rect 10288 32876 10394 32910
rect 10428 32876 10466 32910
rect 10500 32876 10538 32910
rect 10572 32876 10610 32910
rect 10644 32876 10735 32910
rect 10769 32876 10807 32910
rect 10841 32876 10879 32910
rect 10913 32876 10951 32910
rect 10985 32876 11023 32910
rect 11057 32896 11511 32910
rect 11545 32896 11584 32930
rect 11618 32896 11657 32930
rect 11691 32896 11729 32930
rect 11763 32896 11801 32930
rect 11835 32896 11873 32930
rect 11907 32896 11945 32930
rect 11979 32896 11995 32930
rect 11057 32886 11995 32896
rect 12038 32939 15647 32940
rect 12038 32930 13374 32939
rect 13426 32930 13438 32939
rect 13490 32930 13502 32939
rect 12038 32896 12067 32930
rect 12101 32896 12140 32930
rect 12174 32896 12213 32930
rect 12247 32896 12285 32930
rect 12319 32896 12357 32930
rect 12391 32896 12429 32930
rect 12463 32896 12501 32930
rect 12535 32896 12623 32930
rect 12657 32896 12695 32930
rect 12729 32896 12767 32930
rect 12801 32896 12839 32930
rect 12873 32896 12911 32930
rect 12945 32896 12984 32930
rect 13018 32896 13057 32930
rect 13091 32896 13285 32930
rect 13319 32896 13357 32930
rect 13426 32896 13429 32930
rect 13490 32896 13501 32930
rect 12038 32887 13374 32896
rect 13426 32887 13438 32896
rect 13490 32887 13502 32896
rect 13554 32887 13566 32939
rect 13618 32887 13630 32939
rect 13682 32887 13694 32939
rect 13746 32930 15647 32939
rect 13753 32896 13841 32930
rect 13875 32896 13914 32930
rect 13948 32896 13987 32930
rect 14021 32896 14059 32930
rect 14093 32896 14131 32930
rect 14165 32896 14203 32930
rect 14237 32896 14275 32930
rect 14309 32896 15647 32930
rect 13746 32887 15647 32896
rect 15799 32890 15910 32944
rect 16140 32890 16376 32936
rect 12038 32886 15647 32887
rect 11057 32876 11328 32886
rect 9623 32866 11328 32876
rect 8179 32765 8283 32819
rect 8738 32766 8800 32820
rect 8734 32764 8826 32766
rect 9050 32764 9402 32820
rect 8870 32718 8938 32726
rect 8870 32666 8878 32718
rect 8930 32666 8938 32718
rect 8870 32656 8938 32666
rect 5612 31858 5782 32280
rect 5836 31856 6006 32278
rect 6058 31858 6224 32280
rect 6282 31858 6452 32280
rect 6508 31858 6678 32280
rect 9522 31838 9550 32766
rect 11070 32586 11140 32590
rect 11070 32534 11080 32586
rect 11132 32534 11140 32586
rect 11070 32530 11140 32534
rect 16500 32452 16762 33122
rect 16824 32454 17086 33124
rect 17148 32454 17410 33125
rect 17472 32454 17734 33125
rect 17796 32452 18058 33123
rect 18120 32454 18382 33125
rect 18444 32452 18706 33123
rect 18768 32454 19030 33125
rect 21836 33062 21855 33312
rect 22249 33062 22268 33312
rect 21836 33046 22268 33062
rect 23356 33312 23788 33328
rect 23356 33062 23374 33312
rect 23768 33062 23788 33312
rect 21836 32982 22268 32996
rect 19228 32428 19814 32850
rect 19876 32430 20462 32852
rect 20524 32430 21110 32852
rect 21172 32430 21496 32852
rect 21836 32732 21855 32982
rect 22249 32732 22268 32982
rect 21836 32650 22268 32732
rect 23356 32982 23788 33062
rect 23356 32732 23374 32982
rect 23768 32732 23788 32982
rect 23356 32716 23788 32732
rect 21836 32400 21855 32650
rect 22249 32400 22268 32650
rect 21836 32384 22268 32400
rect 23356 32650 23788 32668
rect 23356 32400 23374 32650
rect 23768 32400 23788 32650
rect 11168 31996 11196 32352
rect 10002 31968 11196 31996
rect 7192 31712 7501 31814
rect 9522 31810 10714 31838
rect 6662 30896 7366 30922
rect 6662 30716 6733 30896
rect 6913 30850 7366 30896
rect 6913 30796 7919 30850
rect 6913 30716 7366 30796
rect 6662 30686 7366 30716
rect 6662 30684 7364 30686
rect 9522 30506 9550 31810
rect 9646 31482 11115 31684
rect 9674 31346 10330 31356
rect 9674 31312 9690 31346
rect 9724 31312 9768 31346
rect 9802 31312 9846 31346
rect 9880 31312 9924 31346
rect 9958 31312 10046 31346
rect 10080 31312 10124 31346
rect 10158 31312 10202 31346
rect 10236 31312 10280 31346
rect 10314 31312 10330 31346
rect 9674 31302 10330 31312
rect 10386 31346 11042 31356
rect 10386 31312 10402 31346
rect 10436 31312 10480 31346
rect 10514 31312 10558 31346
rect 10592 31312 10636 31346
rect 10670 31312 10758 31346
rect 10792 31312 10836 31346
rect 10870 31312 10914 31346
rect 10948 31312 10992 31346
rect 11026 31312 11042 31346
rect 10386 31302 11042 31312
rect 10687 31265 10741 31302
rect 9974 31211 10741 31265
rect 9974 31172 10028 31211
rect 9674 31162 10330 31172
rect 9674 31128 9690 31162
rect 9724 31128 9768 31162
rect 9802 31128 9846 31162
rect 9880 31128 9924 31162
rect 9958 31128 10046 31162
rect 10080 31128 10124 31162
rect 10158 31128 10202 31162
rect 10236 31128 10280 31162
rect 10314 31128 10330 31162
rect 9674 31118 10330 31128
rect 10386 31162 11042 31172
rect 10386 31128 10402 31162
rect 10436 31128 10480 31162
rect 10514 31128 10558 31162
rect 10592 31128 10636 31162
rect 10670 31128 10758 31162
rect 10792 31128 10836 31162
rect 10870 31128 10914 31162
rect 10948 31128 10992 31162
rect 11026 31128 11042 31162
rect 10386 31118 11042 31128
rect 11087 30992 11115 31482
rect 9595 30790 9623 30992
rect 9646 30790 11115 30992
rect 11168 30660 11196 31968
rect 21836 32322 22268 32338
rect 21836 32072 21855 32322
rect 22249 32072 22268 32322
rect 21836 31992 22268 32072
rect 23356 32322 23788 32400
rect 23356 32072 23374 32322
rect 23768 32072 23788 32322
rect 23356 32056 23788 32072
rect 11444 31712 16118 31722
rect 11444 31678 11491 31712
rect 11525 31678 11563 31712
rect 11597 31678 11635 31712
rect 11669 31678 11707 31712
rect 11741 31678 11779 31712
rect 11813 31678 11851 31712
rect 11885 31678 11923 31712
rect 11957 31678 12051 31712
rect 12085 31678 12123 31712
rect 12157 31678 12195 31712
rect 12229 31678 12267 31712
rect 12301 31678 12339 31712
rect 12373 31678 12411 31712
rect 12445 31678 12483 31712
rect 12517 31678 12592 31712
rect 12626 31678 12664 31712
rect 12698 31678 12736 31712
rect 12770 31678 12808 31712
rect 12842 31678 12880 31712
rect 12914 31678 12952 31712
rect 12986 31678 13024 31712
rect 13058 31678 13096 31712
rect 13130 31678 13246 31712
rect 13280 31678 13318 31712
rect 13352 31678 13390 31712
rect 13424 31678 13462 31712
rect 13496 31678 13534 31712
rect 13568 31678 13606 31712
rect 13640 31678 13678 31712
rect 13712 31678 13750 31712
rect 13784 31678 13863 31712
rect 13897 31678 13935 31712
rect 13969 31678 14007 31712
rect 14041 31678 14079 31712
rect 14113 31678 14151 31712
rect 14185 31678 14223 31712
rect 14257 31678 14295 31712
rect 14329 31678 16118 31712
rect 11444 31668 16118 31678
rect 16182 31721 16254 31732
rect 16182 31669 16190 31721
rect 16242 31669 16254 31721
rect 16182 31662 16254 31669
rect 16500 31516 17088 31938
rect 17148 31516 17736 31938
rect 17794 31516 18382 31938
rect 18444 31516 19032 31938
rect 21836 31742 21855 31992
rect 22249 31742 22268 31992
rect 21836 31726 22268 31742
rect 23356 31992 23788 32008
rect 23356 31742 23374 31992
rect 23768 31742 23788 31992
rect 21836 31662 22268 31678
rect 21836 31412 21855 31662
rect 22249 31412 22268 31662
rect 16430 31335 16864 31356
rect 16430 31250 16459 31335
rect 11854 31240 13230 31250
rect 11376 31197 11446 31206
rect 11376 31145 11385 31197
rect 11437 31145 11446 31197
rect 11854 31188 12556 31240
rect 12608 31232 13230 31240
rect 12608 31198 12817 31232
rect 12851 31198 12889 31232
rect 12923 31198 12961 31232
rect 12995 31198 13033 31232
rect 13067 31198 13105 31232
rect 13139 31198 13177 31232
rect 13211 31198 13230 31232
rect 12608 31188 13230 31198
rect 11854 31180 13230 31188
rect 14058 31232 16459 31250
rect 14058 31198 14076 31232
rect 14110 31198 14148 31232
rect 14182 31198 14220 31232
rect 14254 31198 14292 31232
rect 14326 31198 14364 31232
rect 14398 31198 14436 31232
rect 14470 31198 16459 31232
rect 14058 31180 16459 31198
rect 11376 31138 11446 31145
rect 11522 31132 11722 31148
rect 11522 31080 11605 31132
rect 11657 31080 11722 31132
rect 11522 31066 11722 31080
rect 16430 31091 16459 31180
rect 16831 31091 16864 31335
rect 16430 31072 16864 31091
rect 21836 31332 22268 31412
rect 23356 31662 23788 31742
rect 23356 31412 23374 31662
rect 23768 31412 23788 31662
rect 23356 31396 23788 31412
rect 21836 31082 21855 31332
rect 22249 31082 22268 31332
rect 21836 31066 22268 31082
rect 23361 31332 23782 31338
rect 23361 31082 23374 31332
rect 23768 31082 23782 31332
rect 23361 31076 23782 31082
rect 10714 30632 11196 30660
rect 9522 30478 10002 30506
rect 11486 30488 12098 30920
rect 12996 30488 13608 30920
rect 9974 30200 10030 30202
rect 9974 30138 10048 30200
rect 9974 30104 9985 30138
rect 10019 30131 10048 30138
rect 9974 30079 9986 30104
rect 10038 30079 10048 30131
rect 9974 30067 10048 30079
rect 9974 30066 9986 30067
rect 9974 30032 9985 30066
rect 9974 30015 9986 30032
rect 10038 30015 10048 30067
rect 9974 30003 10048 30015
rect 9974 29994 9986 30003
rect 9974 29960 9985 29994
rect 9974 29951 9986 29960
rect 10038 29951 10048 30003
rect 9974 29939 10048 29951
rect 9974 29922 9986 29939
rect 9974 29888 9985 29922
rect 9974 29887 9986 29888
rect 10038 29887 10048 29939
rect 9974 29875 10048 29887
rect 9974 29850 9986 29875
rect 9974 29816 9985 29850
rect 10038 29823 10048 29875
rect 10019 29816 10048 29823
rect 9974 29784 10048 29816
rect 9623 29598 11093 29608
rect 9623 29564 9659 29598
rect 9693 29564 9731 29598
rect 9765 29564 9803 29598
rect 9837 29564 9875 29598
rect 9909 29564 9947 29598
rect 9981 29564 10072 29598
rect 10106 29564 10144 29598
rect 10178 29564 10216 29598
rect 10250 29564 10288 29598
rect 10322 29564 10411 29598
rect 10445 29564 10483 29598
rect 10517 29564 10555 29598
rect 10589 29564 10627 29598
rect 10661 29564 10735 29598
rect 10769 29564 10807 29598
rect 10841 29564 10879 29598
rect 10913 29564 10951 29598
rect 10985 29564 11023 29598
rect 11057 29564 11093 29598
rect 9623 29554 11093 29564
rect 9701 29384 11762 29438
rect 11496 29012 11762 29384
rect 11496 28960 11595 29012
rect 11647 28960 11762 29012
rect 7520 27756 10708 28238
rect 7520 27620 10406 27756
rect 7520 25668 8132 27620
rect 10096 27512 10406 27620
rect 10586 27512 10708 27756
rect 9026 26727 9246 26738
rect 9026 26547 9046 26727
rect 9226 26547 9246 26727
rect 9026 26536 9246 26547
rect 10096 25668 10708 27512
rect 11496 27542 11762 28960
rect 12592 29275 12842 29286
rect 12592 28903 12595 29275
rect 12839 28903 12842 29275
rect 12592 28892 12842 28903
rect 12586 28418 13598 28448
rect 12586 28046 12595 28418
rect 12839 28046 13598 28418
rect 12586 28022 13598 28046
rect 12592 27835 12842 27846
rect 11496 26276 11758 27542
rect 12592 27463 12595 27835
rect 12839 27463 12842 27835
rect 12592 27452 12842 27463
rect 11502 26268 11752 26276
rect 11502 25896 11505 26268
rect 11749 25896 11752 26268
rect 11502 25884 11752 25896
rect 11832 26267 12082 26278
rect 11832 25895 11835 26267
rect 12079 25895 12082 26267
rect 11832 25884 12082 25895
rect 13006 25796 13266 26096
rect 13336 25872 13598 28022
rect 7520 25050 10834 25668
rect 11826 25636 13266 25796
rect 11826 25532 12088 25636
rect 13012 25549 13262 25560
rect 13012 25177 13015 25549
rect 13259 25177 13262 25549
rect 13012 25166 13262 25177
rect 11486 20526 12098 20958
rect 12996 20526 13608 20958
rect 11583 19116 17300 19134
rect 25708 19117 25802 19120
rect 25708 19116 25738 19117
rect 11583 19080 25738 19116
rect 17246 19065 25738 19080
rect 25790 19065 25802 19117
rect 17246 19062 25802 19065
rect 20437 19060 20491 19062
rect 25708 19058 25802 19062
rect 13002 17998 15666 18200
rect 7618 17611 7688 17644
rect 7618 17559 7626 17611
rect 7678 17559 7688 17611
rect 7618 17530 7688 17559
rect 7734 17382 7904 17804
rect 7956 17380 8126 17802
rect 8182 17380 8352 17802
rect 8406 17380 8576 17802
rect 8676 17524 9254 17644
rect 9588 17602 9688 17644
rect 9588 17550 9614 17602
rect 9666 17550 9688 17602
rect 9588 17530 9688 17550
rect 9154 17452 9254 17524
rect 9154 17400 9178 17452
rect 9230 17400 9254 17452
rect 9154 17390 9254 17400
rect 9612 16006 9666 17530
rect 12262 17522 16410 17724
rect 18102 17597 19414 17631
rect 21087 17586 22428 17644
rect 12036 16146 12913 16200
rect 13302 16146 14092 16200
rect 14110 16146 15456 16200
rect 16222 16146 16612 16200
rect 17038 16146 17528 16200
rect 18403 16146 19135 16200
rect 14368 16011 14570 16146
rect 18733 16065 18787 16146
rect 19502 15998 19582 16200
rect 19591 16156 19636 16200
rect 19761 16156 20625 16200
rect 19764 16146 20625 16156
rect 21314 16146 22100 16200
rect 22643 16146 22756 16200
rect 21746 16065 21800 16146
rect 18514 15972 19582 15998
rect 18512 15958 19582 15972
rect 14139 15818 14663 15872
rect 11669 15761 11872 15815
rect 12000 15761 13091 15815
rect 13098 15761 13345 15815
rect 13369 15761 13581 15815
rect 15103 15800 17880 15854
rect 18512 15838 18778 15958
rect 18516 15792 18778 15838
rect 11669 15686 11723 15761
rect 13527 15723 13581 15761
rect 14368 15527 14570 15660
rect 14248 15325 14760 15527
rect 17040 15332 18770 15504
rect 18830 15388 19436 15820
rect 19478 15388 20084 15820
rect 20126 15388 20732 15820
rect 20790 15791 21256 15818
rect 23385 15817 23439 16200
rect 23677 16146 25380 16200
rect 20790 15419 20793 15791
rect 21037 15616 21256 15791
rect 21359 15617 23439 15817
rect 21037 15614 21206 15616
rect 21037 15598 21152 15614
rect 21037 15419 21040 15522
rect 20790 15408 21040 15419
rect 21348 15506 21406 15520
rect 21348 15472 21360 15506
rect 21394 15472 21406 15506
rect 10595 15276 10671 15287
rect 10595 15224 10608 15276
rect 10660 15224 10671 15276
rect 10595 15215 10671 15224
rect 10882 15171 10946 15176
rect 9921 15170 11033 15171
rect 9921 15118 10888 15170
rect 10940 15118 11033 15170
rect 9921 15117 11033 15118
rect 10882 15112 10946 15117
rect 11669 15085 11723 15123
rect 13527 15085 13581 15167
rect 11669 15031 11862 15085
rect 11977 15031 12142 15085
rect 12506 15031 12833 15085
rect 13095 15031 13345 15085
rect 13352 15031 13581 15085
rect 9062 14804 9116 15020
rect 10046 15012 10106 15030
rect 17040 15017 17184 15332
rect 18420 15330 18770 15332
rect 21348 15330 21406 15472
rect 9788 14978 10057 15012
rect 10091 14978 10106 15012
rect 9788 14976 10106 14978
rect 9514 14804 9602 14812
rect 9062 14752 9524 14804
rect 9576 14752 9602 14804
rect 9062 14246 9116 14752
rect 9514 14744 9602 14752
rect 9704 14717 9814 14976
rect 10046 14964 10106 14976
rect 14093 14946 14586 15000
rect 15932 14963 17188 15017
rect 21564 14924 22150 15346
rect 22212 14924 22798 15346
rect 22860 14924 23446 15346
rect 23514 15311 23764 15322
rect 23514 15050 23517 15311
rect 23508 14939 23517 15050
rect 23761 15050 23764 15311
rect 23761 14939 23770 15050
rect 11268 14808 11368 14850
rect 11074 14804 11368 14808
rect 11074 14794 11300 14804
rect 11074 14760 11108 14794
rect 11142 14760 11300 14794
rect 11074 14752 11300 14760
rect 11352 14752 11368 14804
rect 11074 14744 11368 14752
rect 9378 14626 9458 14648
rect 9378 14574 9392 14626
rect 9444 14574 9458 14626
rect 9704 14615 9913 14717
rect 11268 14714 11368 14744
rect 23848 14670 24280 15282
rect 25438 15234 25622 15242
rect 25438 15054 25440 15234
rect 25620 15054 25622 15234
rect 25438 15046 25622 15054
rect 9704 14611 9814 14615
rect 9704 14588 9738 14611
rect 9378 14558 9458 14574
rect 10540 14574 10604 14586
rect 10540 14522 10546 14574
rect 10598 14522 10604 14574
rect 13286 14544 13633 14564
rect 10540 14516 10604 14522
rect 11723 14510 13633 14544
rect 14050 14510 17659 14564
rect 17811 14514 17922 14568
rect 18152 14514 18388 14560
rect 11723 14490 13340 14510
rect 10191 14389 10295 14443
rect 10750 14390 10812 14444
rect 10746 14388 10838 14390
rect 11062 14388 11414 14444
rect 10882 14342 10950 14350
rect 10882 14290 10890 14342
rect 10942 14290 10950 14342
rect 10882 14280 10950 14290
rect 7624 13482 7794 13904
rect 7848 13480 8018 13902
rect 8070 13482 8236 13904
rect 8294 13482 8464 13904
rect 8520 13482 8690 13904
rect 11534 13462 11562 14390
rect 13082 14210 13152 14214
rect 13082 14158 13092 14210
rect 13144 14158 13152 14210
rect 13082 14154 13152 14158
rect 13180 13620 13208 13976
rect 18516 13973 18778 14650
rect 18840 13973 19102 14650
rect 19164 13973 19426 14650
rect 19488 13973 19750 14650
rect 19812 13973 20074 14650
rect 20136 13973 20398 14650
rect 20460 13973 20722 14650
rect 20784 13974 21046 14651
rect 21240 14052 21826 14474
rect 21888 14054 22474 14476
rect 22536 14054 23122 14476
rect 23184 14054 23508 14476
rect 23848 14008 24280 14620
rect 25368 14340 25800 14952
rect 12014 13592 13208 13620
rect 9204 13336 9513 13438
rect 11534 13434 12726 13462
rect 7328 12478 9372 12534
rect 7328 12362 7407 12478
rect 7523 12475 9372 12478
rect 7523 12369 9191 12475
rect 9297 12474 9372 12475
rect 9297 12420 9931 12474
rect 9297 12369 9372 12420
rect 7523 12362 9372 12369
rect 7328 12302 9372 12362
rect 11534 12130 11562 13434
rect 11658 13106 13127 13308
rect 11713 12926 11882 12980
rect 11884 12926 12278 12980
rect 12652 12926 12931 12980
rect 12968 12926 13027 12980
rect 12699 12889 12753 12926
rect 11986 12835 12753 12889
rect 11986 12796 12040 12835
rect 11857 12742 12107 12796
rect 12553 12742 12942 12796
rect 13099 12616 13127 13106
rect 11607 12414 11635 12616
rect 11658 12414 13127 12616
rect 13180 12284 13208 13592
rect 18202 13346 18280 13356
rect 13486 13292 18130 13346
rect 18202 13294 18216 13346
rect 18268 13294 18280 13346
rect 18202 13288 18280 13294
rect 18516 13036 19102 13458
rect 19164 13036 19750 13458
rect 19812 13036 20398 13458
rect 20460 13036 21046 13458
rect 23848 13350 24280 13962
rect 25368 13680 25800 14292
rect 18442 12959 18876 12980
rect 18442 12874 18471 12959
rect 13866 12864 15242 12874
rect 13388 12821 13458 12830
rect 13388 12769 13397 12821
rect 13449 12769 13458 12821
rect 13866 12812 14568 12864
rect 14620 12812 15242 12864
rect 13866 12804 15242 12812
rect 16070 12804 18471 12874
rect 13388 12762 13458 12769
rect 13534 12756 13734 12772
rect 13534 12704 13617 12756
rect 13669 12704 13734 12756
rect 13534 12690 13734 12704
rect 18442 12715 18471 12804
rect 18843 12715 18876 12959
rect 18442 12696 18876 12715
rect 23848 12690 24280 13302
rect 25368 13020 25800 13632
rect 25386 12953 25780 12956
rect 25386 12709 25397 12953
rect 25769 12709 25780 12953
rect 25386 12706 25780 12709
rect 12726 12256 13208 12284
rect 11534 12102 12014 12130
rect 13498 12112 14110 12544
rect 15008 12112 15620 12544
rect 11986 11824 12042 11826
rect 11986 11762 12060 11824
rect 11986 11728 11997 11762
rect 12031 11755 12060 11762
rect 11986 11703 11998 11728
rect 12050 11703 12060 11755
rect 11986 11691 12060 11703
rect 11986 11690 11998 11691
rect 11986 11656 11997 11690
rect 11986 11639 11998 11656
rect 12050 11639 12060 11691
rect 11986 11627 12060 11639
rect 11986 11618 11998 11627
rect 11986 11584 11997 11618
rect 11986 11575 11998 11584
rect 12050 11575 12060 11627
rect 11986 11563 12060 11575
rect 11986 11546 11998 11563
rect 11986 11512 11997 11546
rect 11986 11511 11998 11512
rect 12050 11511 12060 11563
rect 11986 11499 12060 11511
rect 11986 11474 11998 11499
rect 11986 11440 11997 11474
rect 12050 11447 12060 11499
rect 12031 11440 12060 11447
rect 11986 11408 12060 11440
rect 11642 11178 13094 11232
rect 11713 11008 13774 11062
rect 13508 10636 13774 11008
rect 13508 10584 13607 10636
rect 13659 10584 13774 10636
rect 9532 9380 12720 9862
rect 9532 9244 12418 9380
rect 9532 7292 10144 9244
rect 12108 9136 12418 9244
rect 12598 9136 12720 9380
rect 11038 8351 11258 8362
rect 11038 8171 11058 8351
rect 11238 8171 11258 8351
rect 11038 8160 11258 8171
rect 12108 7292 12720 9136
rect 13508 9166 13774 10584
rect 14604 10899 14854 10910
rect 14604 10527 14607 10899
rect 14851 10527 14854 10899
rect 14604 10516 14854 10527
rect 14598 10042 15610 10072
rect 14598 9670 14607 10042
rect 14851 9670 15610 10042
rect 14598 9646 15610 9670
rect 14604 9459 14854 9470
rect 13508 7900 13770 9166
rect 14604 9087 14607 9459
rect 14851 9087 14854 9459
rect 14604 9076 14854 9087
rect 13514 7892 13764 7900
rect 13514 7520 13517 7892
rect 13761 7520 13764 7892
rect 13514 7508 13764 7520
rect 13844 7891 14094 7902
rect 13844 7519 13847 7891
rect 14091 7519 14094 7891
rect 13844 7508 14094 7519
rect 15018 7420 15278 7720
rect 15348 7496 15610 9646
rect 9532 6674 12846 7292
rect 13838 7260 15278 7420
rect 13838 7156 14100 7260
rect 15024 7173 15274 7184
rect 15024 6801 15027 7173
rect 15271 6801 15274 7173
rect 15024 6790 15274 6801
rect 13498 2150 14110 2582
rect 15008 2150 15620 2582
<< via1 >>
rect 5614 35935 5666 35987
rect 7602 35926 7654 35978
rect 7166 35776 7218 35828
rect 9029 34357 9081 34409
rect 8596 33644 8648 33654
rect 8596 33610 8606 33644
rect 8606 33610 8640 33644
rect 8640 33610 8648 33644
rect 8596 33602 8648 33610
rect 8870 33493 8922 33545
rect 18777 33889 19021 34261
rect 7512 33172 7564 33180
rect 7512 33138 7521 33172
rect 7521 33138 7555 33172
rect 7555 33138 7564 33172
rect 7512 33128 7564 33138
rect 21505 33315 21749 33687
rect 23428 33430 23608 33610
rect 23670 33556 23722 33608
rect 23670 33486 23722 33538
rect 23670 33416 23722 33468
rect 9288 33128 9340 33180
rect 7380 32993 7432 33002
rect 7380 32959 7389 32993
rect 7389 32959 7423 32993
rect 7423 32959 7432 32993
rect 7380 32950 7432 32959
rect 8534 32946 8586 32950
rect 8534 32912 8542 32946
rect 8542 32912 8576 32946
rect 8576 32912 8586 32946
rect 8534 32898 8586 32912
rect 13374 32930 13426 32939
rect 13438 32930 13490 32939
rect 13502 32930 13554 32939
rect 13374 32896 13391 32930
rect 13391 32896 13426 32930
rect 13438 32896 13463 32930
rect 13463 32896 13490 32930
rect 13502 32896 13535 32930
rect 13535 32896 13554 32930
rect 13374 32887 13426 32896
rect 13438 32887 13490 32896
rect 13502 32887 13554 32896
rect 13566 32930 13618 32939
rect 13566 32896 13573 32930
rect 13573 32896 13607 32930
rect 13607 32896 13618 32930
rect 13566 32887 13618 32896
rect 13630 32930 13682 32939
rect 13630 32896 13646 32930
rect 13646 32896 13680 32930
rect 13680 32896 13682 32930
rect 13630 32887 13682 32896
rect 13694 32930 13746 32939
rect 13694 32896 13719 32930
rect 13719 32896 13746 32930
rect 13694 32887 13746 32896
rect 8878 32710 8930 32718
rect 8878 32676 8886 32710
rect 8886 32676 8920 32710
rect 8920 32676 8930 32710
rect 8878 32666 8930 32676
rect 11080 32578 11132 32586
rect 11080 32544 11091 32578
rect 11091 32544 11125 32578
rect 11125 32544 11132 32578
rect 11080 32534 11132 32544
rect 6733 30716 6913 30896
rect 16190 31669 16242 31721
rect 11385 31190 11437 31197
rect 11385 31156 11396 31190
rect 11396 31156 11430 31190
rect 11430 31156 11437 31190
rect 11385 31145 11437 31156
rect 12556 31188 12608 31240
rect 11605 31080 11657 31132
rect 16459 31091 16831 31335
rect 23385 31085 23757 31329
rect 9986 30104 10019 30131
rect 10019 30104 10038 30131
rect 9986 30079 10038 30104
rect 9986 30066 10038 30067
rect 9986 30032 10019 30066
rect 10019 30032 10038 30066
rect 9986 30015 10038 30032
rect 9986 29994 10038 30003
rect 9986 29960 10019 29994
rect 10019 29960 10038 29994
rect 9986 29951 10038 29960
rect 9986 29922 10038 29939
rect 9986 29888 10019 29922
rect 10019 29888 10038 29922
rect 9986 29887 10038 29888
rect 9986 29850 10038 29875
rect 9986 29823 10019 29850
rect 10019 29823 10038 29850
rect 11595 28960 11647 29012
rect 10406 27512 10586 27756
rect 9046 26547 9226 26727
rect 12595 28046 12839 28418
rect 12595 27463 12839 27835
rect 11505 25896 11749 26268
rect 11835 25895 12079 26267
rect 13015 25177 13259 25549
rect 25738 19065 25790 19117
rect 7626 17559 7678 17611
rect 9614 17550 9666 17602
rect 9178 17400 9230 17452
rect 20793 15419 21037 15791
rect 10608 15268 10660 15276
rect 10608 15234 10618 15268
rect 10618 15234 10652 15268
rect 10652 15234 10660 15268
rect 10608 15224 10660 15234
rect 10888 15118 10940 15170
rect 9524 14796 9576 14804
rect 9524 14762 9533 14796
rect 9533 14762 9567 14796
rect 9567 14762 9576 14796
rect 9524 14752 9576 14762
rect 23517 14939 23761 15311
rect 11300 14752 11352 14804
rect 9392 14617 9444 14626
rect 9392 14583 9401 14617
rect 9401 14583 9435 14617
rect 9435 14583 9444 14617
rect 9392 14574 9444 14583
rect 25440 15054 25620 15234
rect 25682 15180 25734 15232
rect 25682 15110 25734 15162
rect 25682 15040 25734 15092
rect 10546 14570 10598 14574
rect 10546 14536 10554 14570
rect 10554 14536 10588 14570
rect 10588 14536 10598 14570
rect 10546 14522 10598 14536
rect 10890 14334 10942 14342
rect 10890 14300 10898 14334
rect 10898 14300 10932 14334
rect 10932 14300 10942 14334
rect 10890 14290 10942 14300
rect 13092 14202 13144 14210
rect 13092 14168 13103 14202
rect 13103 14168 13137 14202
rect 13137 14168 13144 14202
rect 13092 14158 13144 14168
rect 7407 12362 7523 12478
rect 18216 13294 18268 13346
rect 13397 12814 13449 12821
rect 13397 12780 13408 12814
rect 13408 12780 13442 12814
rect 13442 12780 13449 12814
rect 13397 12769 13449 12780
rect 14568 12812 14620 12864
rect 13617 12704 13669 12756
rect 18471 12715 18843 12959
rect 25397 12709 25769 12953
rect 11998 11728 12031 11755
rect 12031 11728 12050 11755
rect 11998 11703 12050 11728
rect 11998 11690 12050 11691
rect 11998 11656 12031 11690
rect 12031 11656 12050 11690
rect 11998 11639 12050 11656
rect 11998 11618 12050 11627
rect 11998 11584 12031 11618
rect 12031 11584 12050 11618
rect 11998 11575 12050 11584
rect 11998 11546 12050 11563
rect 11998 11512 12031 11546
rect 12031 11512 12050 11546
rect 11998 11511 12050 11512
rect 11998 11474 12050 11499
rect 11998 11447 12031 11474
rect 12031 11447 12050 11474
rect 13607 10584 13659 10636
rect 12418 9136 12598 9380
rect 11058 8171 11238 8351
rect 14607 9670 14851 10042
rect 14607 9087 14851 9459
rect 13517 7520 13761 7892
rect 13847 7519 14091 7891
rect 15027 6801 15271 7173
<< metal2 >>
rect 5596 35987 7676 36020
rect 5596 35935 5614 35987
rect 5666 35978 7676 35987
rect 5666 35935 7602 35978
rect 5596 35926 7602 35935
rect 7654 35926 7676 35978
rect 15436 35973 18058 36007
rect 18448 35975 23696 36009
rect 5596 35906 7676 35926
rect 7142 35828 7242 35846
rect 7142 35776 7166 35828
rect 7218 35776 7242 35828
rect 7142 32922 7242 35776
rect 10901 34522 13822 34576
rect 15916 34522 17579 34576
rect 18906 34522 20631 34576
rect 9006 34412 9102 34456
rect 12356 34414 19761 34468
rect 9006 34356 9026 34412
rect 9082 34356 9102 34412
rect 9006 34312 9102 34356
rect 12356 34036 12558 34387
rect 18766 34261 19030 34284
rect 18766 33889 18777 34261
rect 19021 33889 19030 34261
rect 8568 33654 8672 33678
rect 8568 33598 8592 33654
rect 8648 33598 8672 33654
rect 8568 33576 8672 33598
rect 8848 33547 8944 33568
rect 10652 33562 10680 33628
rect 8848 33491 8868 33547
rect 8924 33491 8944 33547
rect 8848 33470 8944 33491
rect 9522 33534 12117 33562
rect 7486 33182 7590 33204
rect 7486 33126 7510 33182
rect 7566 33126 7590 33182
rect 7486 33104 7590 33126
rect 9256 33182 9356 33226
rect 9256 33126 9286 33182
rect 9342 33126 9356 33182
rect 9256 33090 9356 33126
rect 7366 33004 7446 33024
rect 7366 32948 7378 33004
rect 7434 32948 7446 33004
rect 7366 32934 7446 32948
rect 8528 32950 8592 32962
rect 8528 32898 8534 32950
rect 8586 32898 8592 32950
rect 8528 32892 8592 32898
rect 8534 32726 8586 32892
rect 9522 32769 9550 33534
rect 11156 33447 11196 33448
rect 10794 33419 11196 33447
rect 11140 33418 11196 33419
rect 8534 32718 8938 32726
rect 8534 32666 8878 32718
rect 8930 32666 8938 32718
rect 8534 32656 8938 32666
rect 6660 30896 6976 30922
rect 6660 30875 6733 30896
rect 6913 30875 6976 30896
rect 6660 30739 6713 30875
rect 6929 30739 6976 30875
rect 6660 30716 6733 30739
rect 6913 30716 6976 30739
rect 6660 30684 6976 30716
rect 9674 29411 9728 33117
rect 9974 31265 10028 31329
rect 9974 31211 10749 31265
rect 10695 31145 10749 31211
rect 9974 30131 10048 30202
rect 9974 30125 9986 30131
rect 10038 30125 10048 30131
rect 9974 30069 9984 30125
rect 10040 30069 10048 30125
rect 9974 30067 10048 30069
rect 9974 30045 9986 30067
rect 10038 30045 10048 30067
rect 9974 29989 9984 30045
rect 10040 29989 10048 30045
rect 9974 29965 9986 29989
rect 10038 29965 10048 29989
rect 9974 29909 9984 29965
rect 10040 29909 10048 29965
rect 9974 29887 9986 29909
rect 10038 29887 10048 29909
rect 9974 29885 10048 29887
rect 9974 29829 9984 29885
rect 10040 29829 10048 29885
rect 9974 29823 9986 29829
rect 10038 29823 10048 29829
rect 9974 29784 10048 29823
rect 10988 29496 11042 33119
rect 11070 32590 11134 32600
rect 11070 32534 11078 32590
rect 11070 32524 11134 32534
rect 11168 32346 11196 33418
rect 12089 33349 12117 33534
rect 12547 32339 12611 33802
rect 13875 32939 13909 33847
rect 18766 33712 19030 33889
rect 18766 33687 21758 33712
rect 18766 33315 21505 33687
rect 21749 33315 21758 33687
rect 23556 33658 23722 35276
rect 23356 33610 23788 33658
rect 23356 33430 23428 33610
rect 23608 33608 23788 33610
rect 23608 33556 23670 33608
rect 23722 33556 23788 33608
rect 23608 33538 23788 33556
rect 23608 33486 23670 33538
rect 23722 33486 23788 33538
rect 23608 33468 23788 33486
rect 23608 33430 23670 33468
rect 23356 33416 23670 33430
rect 23722 33416 23788 33468
rect 23356 33376 23788 33416
rect 18766 33286 21758 33315
rect 13368 32887 13374 32939
rect 13426 32887 13438 32939
rect 13490 32887 13502 32939
rect 13554 32887 13566 32939
rect 13618 32887 13630 32939
rect 13682 32887 13694 32939
rect 13746 32887 14135 32939
rect 12547 32305 15119 32339
rect 12547 31250 12611 32305
rect 21496 31740 21758 33286
rect 16170 31721 21758 31740
rect 16170 31669 16190 31721
rect 16242 31669 21758 31721
rect 16170 31650 21758 31669
rect 16430 31335 16864 31356
rect 16430 31321 16459 31335
rect 16831 31321 16864 31335
rect 12546 31240 12612 31250
rect 11372 31199 11450 31210
rect 11372 31143 11383 31199
rect 11439 31143 11450 31199
rect 12546 31188 12556 31240
rect 12608 31188 12612 31240
rect 12546 31180 12612 31188
rect 11372 31134 11450 31143
rect 11522 31134 11722 31148
rect 11522 31078 11603 31134
rect 11659 31078 11722 31134
rect 11522 31066 11722 31078
rect 16430 31105 16457 31321
rect 16833 31105 16864 31321
rect 16430 31091 16459 31105
rect 16831 31091 16864 31105
rect 16430 31072 16864 31091
rect 21496 31338 21758 31650
rect 21496 31329 23782 31338
rect 21496 31085 23385 31329
rect 23757 31085 23782 31329
rect 21496 31076 23782 31085
rect 10988 29436 12850 29496
rect 11522 29014 11722 29052
rect 11522 28958 11593 29014
rect 11649 28958 11722 29014
rect 11522 28916 11722 28958
rect 12586 28418 12850 29436
rect 12586 28046 12595 28418
rect 12839 28046 12850 28418
rect 12586 28022 12850 28046
rect 10294 27835 12848 27860
rect 10294 27756 12595 27835
rect 10294 27512 10406 27756
rect 10586 27512 12595 27756
rect 10294 27463 12595 27512
rect 12839 27463 12848 27835
rect 10294 27438 12848 27463
rect 8986 26727 11758 26756
rect 8986 26547 9046 26727
rect 9226 26547 11758 26727
rect 8986 26510 11758 26547
rect 11496 26268 11758 26510
rect 11496 25896 11505 26268
rect 11749 25896 11758 26268
rect 11496 25870 11758 25896
rect 11826 26267 12088 26292
rect 11826 25895 11835 26267
rect 12079 25895 12088 26267
rect 11826 25872 12088 25895
rect 11826 25796 12086 25872
rect 11826 25636 13266 25796
rect 13006 25574 13266 25636
rect 13006 25549 13268 25574
rect 13006 25177 13015 25549
rect 13259 25177 13268 25549
rect 13006 25154 13268 25177
rect 25716 19117 25812 19134
rect 25716 19116 25738 19117
rect 25790 19116 25812 19117
rect 25716 19060 25736 19116
rect 25792 19060 25812 19116
rect 25716 19042 25812 19060
rect 7608 17611 9688 17644
rect 7608 17559 7626 17611
rect 7678 17602 9688 17611
rect 7678 17559 9614 17602
rect 7608 17550 9614 17559
rect 9666 17550 9688 17602
rect 17448 17597 20070 17631
rect 20460 17599 25708 17633
rect 7608 17530 9688 17550
rect 9154 17452 9254 17470
rect 9154 17400 9178 17452
rect 9230 17400 9254 17452
rect 9154 14546 9254 17400
rect 12913 16146 15834 16200
rect 17928 16146 19591 16200
rect 20918 16146 22643 16200
rect 14368 16038 21773 16092
rect 14368 15660 14570 16011
rect 20782 15791 21046 15814
rect 10590 15278 10676 15296
rect 10590 15222 10606 15278
rect 10662 15222 10676 15278
rect 10590 15206 10676 15222
rect 10862 15172 10966 15196
rect 12664 15186 12692 15252
rect 10862 15116 10885 15172
rect 10941 15116 10966 15172
rect 10862 15092 10966 15116
rect 11534 15158 14129 15186
rect 9500 14806 9598 14826
rect 9500 14750 9521 14806
rect 9577 14750 9598 14806
rect 9500 14730 9598 14750
rect 11268 14806 11368 14850
rect 11268 14750 11298 14806
rect 11354 14750 11368 14806
rect 11268 14714 11368 14750
rect 9378 14628 9458 14648
rect 9378 14572 9390 14628
rect 9446 14572 9458 14628
rect 9378 14558 9458 14572
rect 10540 14574 10604 14586
rect 10540 14522 10546 14574
rect 10598 14522 10604 14574
rect 10540 14516 10604 14522
rect 10546 14350 10598 14516
rect 11534 14393 11562 15158
rect 13168 15071 13208 15072
rect 12806 15043 13208 15071
rect 13152 15042 13208 15043
rect 10546 14342 10950 14350
rect 10546 14290 10890 14342
rect 10942 14290 10950 14342
rect 10546 14280 10950 14290
rect 7374 12489 7552 12508
rect 7374 12353 7396 12489
rect 7532 12353 7552 12489
rect 7374 12330 7552 12353
rect 11686 11035 11740 14741
rect 11986 12889 12040 12953
rect 11986 12835 12761 12889
rect 12707 12769 12761 12835
rect 11986 11755 12060 11826
rect 11986 11749 11998 11755
rect 12050 11749 12060 11755
rect 11986 11693 11996 11749
rect 12052 11693 12060 11749
rect 11986 11691 12060 11693
rect 11986 11669 11998 11691
rect 12050 11669 12060 11691
rect 11986 11613 11996 11669
rect 12052 11613 12060 11669
rect 11986 11589 11998 11613
rect 12050 11589 12060 11613
rect 11986 11533 11996 11589
rect 12052 11533 12060 11589
rect 11986 11511 11998 11533
rect 12050 11511 12060 11533
rect 11986 11509 12060 11511
rect 11986 11453 11996 11509
rect 12052 11453 12060 11509
rect 11986 11447 11998 11453
rect 12050 11447 12060 11453
rect 11986 11408 12060 11447
rect 13000 11120 13054 14743
rect 13082 14214 13146 14224
rect 13082 14158 13090 14214
rect 13082 14148 13146 14158
rect 13180 13970 13208 15042
rect 14101 14973 14129 15158
rect 14559 13963 14623 15426
rect 15887 14563 15921 15471
rect 20782 15419 20793 15791
rect 21037 15419 21046 15791
rect 20782 15336 21046 15419
rect 20782 15311 23770 15336
rect 20782 14939 23517 15311
rect 23761 14939 23770 15311
rect 25568 15282 25734 16900
rect 25368 15234 25800 15282
rect 25368 15054 25440 15234
rect 25620 15232 25800 15234
rect 25620 15180 25682 15232
rect 25734 15180 25800 15232
rect 25620 15162 25800 15180
rect 25620 15110 25682 15162
rect 25734 15110 25800 15162
rect 25620 15092 25800 15110
rect 25620 15054 25682 15092
rect 25368 15040 25682 15054
rect 25734 15040 25800 15092
rect 25368 15000 25800 15040
rect 20782 14910 23770 14939
rect 15572 14511 16147 14563
rect 14559 13929 17131 13963
rect 14559 12874 14623 13929
rect 23508 13356 23770 14910
rect 18202 13346 23770 13356
rect 18202 13294 18216 13346
rect 18268 13294 23770 13346
rect 18202 13288 23770 13294
rect 18442 12959 18876 12980
rect 18442 12945 18471 12959
rect 18843 12945 18876 12959
rect 14558 12864 14624 12874
rect 13384 12823 13462 12834
rect 13384 12767 13395 12823
rect 13451 12767 13462 12823
rect 14558 12812 14568 12864
rect 14620 12812 14624 12864
rect 14558 12804 14624 12812
rect 13384 12758 13462 12767
rect 13534 12758 13734 12772
rect 13534 12702 13615 12758
rect 13671 12702 13734 12758
rect 13534 12690 13734 12702
rect 18442 12729 18469 12945
rect 18845 12729 18876 12945
rect 18442 12715 18471 12729
rect 18843 12715 18876 12729
rect 18442 12696 18876 12715
rect 23508 12962 23770 13288
rect 23508 12953 25794 12962
rect 23508 12709 25397 12953
rect 25769 12709 25794 12953
rect 23508 12700 25794 12709
rect 13000 11060 14862 11120
rect 13534 10638 13734 10676
rect 13534 10582 13605 10638
rect 13661 10582 13734 10638
rect 13534 10540 13734 10582
rect 14598 10042 14862 11060
rect 14598 9670 14607 10042
rect 14851 9670 14862 10042
rect 14598 9646 14862 9670
rect 12306 9459 14860 9484
rect 12306 9380 14607 9459
rect 12306 9136 12418 9380
rect 12598 9136 14607 9380
rect 12306 9087 14607 9136
rect 14851 9087 14860 9459
rect 12306 9062 14860 9087
rect 10998 8351 13770 8380
rect 10998 8171 11058 8351
rect 11238 8171 13770 8351
rect 10998 8134 13770 8171
rect 13508 7892 13770 8134
rect 13508 7520 13517 7892
rect 13761 7520 13770 7892
rect 13508 7494 13770 7520
rect 13838 7891 14100 7916
rect 13838 7519 13847 7891
rect 14091 7519 14100 7891
rect 13838 7496 14100 7519
rect 13838 7420 14098 7496
rect 13838 7260 15278 7420
rect 15018 7198 15278 7260
rect 15018 7173 15280 7198
rect 15018 6801 15027 7173
rect 15271 6801 15280 7173
rect 15018 6778 15280 6801
<< via2 >>
rect 9026 34409 9082 34412
rect 9026 34357 9029 34409
rect 9029 34357 9081 34409
rect 9081 34357 9082 34409
rect 9026 34356 9082 34357
rect 8592 33602 8596 33654
rect 8596 33602 8648 33654
rect 8592 33598 8648 33602
rect 8868 33545 8924 33547
rect 8868 33493 8870 33545
rect 8870 33493 8922 33545
rect 8922 33493 8924 33545
rect 8868 33491 8924 33493
rect 7510 33180 7566 33182
rect 7510 33128 7512 33180
rect 7512 33128 7564 33180
rect 7564 33128 7566 33180
rect 7510 33126 7566 33128
rect 9286 33180 9342 33182
rect 9286 33128 9288 33180
rect 9288 33128 9340 33180
rect 9340 33128 9342 33180
rect 9286 33126 9342 33128
rect 7378 33002 7434 33004
rect 7378 32950 7380 33002
rect 7380 32950 7432 33002
rect 7432 32950 7434 33002
rect 7378 32948 7434 32950
rect 6713 30739 6733 30875
rect 6733 30739 6913 30875
rect 6913 30739 6929 30875
rect 9984 30079 9986 30125
rect 9986 30079 10038 30125
rect 10038 30079 10040 30125
rect 9984 30069 10040 30079
rect 9984 30015 9986 30045
rect 9986 30015 10038 30045
rect 10038 30015 10040 30045
rect 9984 30003 10040 30015
rect 9984 29989 9986 30003
rect 9986 29989 10038 30003
rect 10038 29989 10040 30003
rect 9984 29951 9986 29965
rect 9986 29951 10038 29965
rect 10038 29951 10040 29965
rect 9984 29939 10040 29951
rect 9984 29909 9986 29939
rect 9986 29909 10038 29939
rect 10038 29909 10040 29939
rect 9984 29875 10040 29885
rect 9984 29829 9986 29875
rect 9986 29829 10038 29875
rect 10038 29829 10040 29875
rect 11078 32586 11134 32590
rect 11078 32534 11080 32586
rect 11080 32534 11132 32586
rect 11132 32534 11134 32586
rect 23450 33452 23586 33588
rect 11383 31197 11439 31199
rect 11383 31145 11385 31197
rect 11385 31145 11437 31197
rect 11437 31145 11439 31197
rect 11383 31143 11439 31145
rect 11603 31132 11659 31134
rect 11603 31080 11605 31132
rect 11605 31080 11657 31132
rect 11657 31080 11659 31132
rect 11603 31078 11659 31080
rect 16457 31105 16459 31321
rect 16459 31105 16831 31321
rect 16831 31105 16833 31321
rect 11593 29012 11649 29014
rect 11593 28960 11595 29012
rect 11595 28960 11647 29012
rect 11647 28960 11649 29012
rect 11593 28958 11649 28960
rect 25736 19065 25738 19116
rect 25738 19065 25790 19116
rect 25790 19065 25792 19116
rect 25736 19060 25792 19065
rect 10606 15276 10662 15278
rect 10606 15224 10608 15276
rect 10608 15224 10660 15276
rect 10660 15224 10662 15276
rect 10606 15222 10662 15224
rect 10885 15170 10941 15172
rect 10885 15118 10888 15170
rect 10888 15118 10940 15170
rect 10940 15118 10941 15170
rect 10885 15116 10941 15118
rect 9521 14804 9577 14806
rect 9521 14752 9524 14804
rect 9524 14752 9576 14804
rect 9576 14752 9577 14804
rect 9521 14750 9577 14752
rect 11298 14804 11354 14806
rect 11298 14752 11300 14804
rect 11300 14752 11352 14804
rect 11352 14752 11354 14804
rect 11298 14750 11354 14752
rect 9390 14626 9446 14628
rect 9390 14574 9392 14626
rect 9392 14574 9444 14626
rect 9444 14574 9446 14626
rect 9390 14572 9446 14574
rect 7396 12478 7532 12489
rect 7396 12362 7407 12478
rect 7407 12362 7523 12478
rect 7523 12362 7532 12478
rect 7396 12353 7532 12362
rect 11996 11703 11998 11749
rect 11998 11703 12050 11749
rect 12050 11703 12052 11749
rect 11996 11693 12052 11703
rect 11996 11639 11998 11669
rect 11998 11639 12050 11669
rect 12050 11639 12052 11669
rect 11996 11627 12052 11639
rect 11996 11613 11998 11627
rect 11998 11613 12050 11627
rect 12050 11613 12052 11627
rect 11996 11575 11998 11589
rect 11998 11575 12050 11589
rect 12050 11575 12052 11589
rect 11996 11563 12052 11575
rect 11996 11533 11998 11563
rect 11998 11533 12050 11563
rect 12050 11533 12052 11563
rect 11996 11499 12052 11509
rect 11996 11453 11998 11499
rect 11998 11453 12050 11499
rect 12050 11453 12052 11499
rect 13090 14210 13146 14214
rect 13090 14158 13092 14210
rect 13092 14158 13144 14210
rect 13144 14158 13146 14210
rect 25462 15076 25598 15212
rect 13395 12821 13451 12823
rect 13395 12769 13397 12821
rect 13397 12769 13449 12821
rect 13449 12769 13451 12821
rect 13395 12767 13451 12769
rect 13615 12756 13671 12758
rect 13615 12704 13617 12756
rect 13617 12704 13669 12756
rect 13669 12704 13671 12756
rect 13615 12702 13671 12704
rect 18469 12729 18471 12945
rect 18471 12729 18843 12945
rect 18843 12729 18845 12945
rect 13605 10636 13661 10638
rect 13605 10584 13607 10636
rect 13607 10584 13659 10636
rect 13659 10584 13661 10636
rect 13605 10582 13661 10584
<< metal3 >>
rect 8568 38434 8670 38464
rect 8568 38429 8672 38434
rect 8568 38365 8583 38429
rect 8647 38365 8672 38429
rect 8568 33654 8672 38365
rect 9561 35319 9731 35322
rect 9561 35259 15071 35319
rect 9561 35210 9731 35259
rect 8568 33598 8592 33654
rect 8648 33598 8672 33654
rect 8568 33576 8672 33598
rect 9008 34412 9158 34510
rect 9008 34356 9026 34412
rect 9082 34356 9158 34412
rect 8846 33547 8946 33568
rect 8846 33491 8868 33547
rect 8924 33491 8946 33547
rect 8846 33478 8946 33491
rect 5022 33468 8946 33478
rect 5022 33404 5107 33468
rect 5171 33404 5187 33468
rect 5251 33404 5267 33468
rect 5331 33404 8946 33468
rect 5022 33394 8946 33404
rect 7480 33186 7596 33210
rect 7480 33122 7506 33186
rect 7570 33122 7596 33186
rect 7480 33098 7596 33122
rect 7356 33008 7456 33038
rect 7356 32944 7376 33008
rect 7440 32944 7456 33008
rect 7356 32922 7456 32944
rect 9008 31676 9158 34356
rect 9008 31612 9055 31676
rect 9119 31612 9158 31676
rect 9008 31602 9158 31612
rect 9256 33182 9356 33226
rect 9256 33126 9286 33182
rect 9342 33126 9356 33182
rect 9256 31210 9356 33126
rect 9671 33117 9731 35210
rect 10356 34948 14314 35008
rect 10985 33119 11045 34948
rect 18028 34321 18088 34669
rect 18028 34261 19366 34321
rect 23356 33592 23788 33658
rect 23356 33448 23446 33592
rect 23590 33448 23788 33592
rect 23356 33376 23788 33448
rect 11064 32590 11146 32600
rect 11064 32534 11078 32590
rect 11134 32534 15013 32590
rect 11064 32530 15013 32534
rect 11064 32524 11146 32530
rect 16430 31324 16864 31356
rect 16430 31321 16494 31324
rect 16798 31321 16864 31324
rect 9256 31199 11450 31210
rect 9256 31143 11383 31199
rect 11439 31143 11450 31199
rect 9256 31134 11450 31143
rect 11522 31134 11722 31148
rect 11522 31078 11603 31134
rect 11659 31078 11722 31134
rect 800 30875 6976 30922
rect 800 30874 6713 30875
rect 800 30730 849 30874
rect 993 30739 6713 30874
rect 6929 30739 6976 30875
rect 993 30730 6976 30739
rect 800 30686 6976 30730
rect 800 30682 2806 30686
rect 9974 30132 10060 30202
rect 9974 30125 9988 30132
rect 9974 30069 9984 30125
rect 9974 30068 9988 30069
rect 10052 30068 10060 30132
rect 9974 30045 10060 30068
rect 9974 29989 9984 30045
rect 10040 30030 10060 30045
rect 9974 29966 9990 29989
rect 10054 29966 10060 30030
rect 9974 29965 10060 29966
rect 9974 29909 9984 29965
rect 10040 29918 10060 29965
rect 9974 29885 9988 29909
rect 9974 29829 9984 29885
rect 10052 29854 10060 29918
rect 10040 29829 10060 29854
rect 9974 29784 10060 29829
rect 11522 29014 11722 31078
rect 16430 31105 16457 31321
rect 16833 31105 16864 31321
rect 16430 31100 16494 31105
rect 16798 31100 16864 31105
rect 16430 31072 16864 31100
rect 16430 31070 16833 31072
rect 11522 28958 11593 29014
rect 11649 28958 11722 29014
rect 11522 28916 11722 28958
rect 10582 19966 10686 19988
rect 10582 19902 10602 19966
rect 10666 19902 10686 19966
rect 10582 19884 10686 19902
rect 10584 15282 10682 19884
rect 25714 19120 25814 19136
rect 25714 19056 25732 19120
rect 25796 19056 25814 19120
rect 25714 19038 25814 19056
rect 11573 16943 11743 16946
rect 11573 16883 17083 16943
rect 11573 16834 11743 16883
rect 10584 15218 10602 15282
rect 10666 15218 10682 15282
rect 10584 15202 10682 15218
rect 10862 15172 10966 15196
rect 10862 15116 10885 15172
rect 10941 15116 10966 15172
rect 9496 14810 9602 14830
rect 9496 14746 9517 14810
rect 9581 14746 9602 14810
rect 9496 14726 9602 14746
rect 9368 14632 9468 14662
rect 9368 14568 9388 14632
rect 9452 14568 9468 14632
rect 9368 14546 9468 14568
rect 10862 13796 10966 15116
rect 10862 13732 10882 13796
rect 10946 13732 10966 13796
rect 10862 13700 10966 13732
rect 11268 14806 11368 14850
rect 11268 14750 11298 14806
rect 11354 14750 11368 14806
rect 11268 12834 11368 14750
rect 11683 14741 11743 16834
rect 12368 16572 16326 16632
rect 12997 14743 13057 16572
rect 20040 15945 20100 16293
rect 20040 15885 21378 15945
rect 25368 15216 25800 15282
rect 25368 15072 25458 15216
rect 25602 15072 25800 15216
rect 25368 15000 25800 15072
rect 13076 14214 13158 14224
rect 13076 14158 13090 14214
rect 13146 14158 17025 14214
rect 13076 14154 17025 14158
rect 13076 14148 13158 14154
rect 18442 12948 18876 12980
rect 18442 12945 18506 12948
rect 18810 12945 18876 12948
rect 11268 12823 13462 12834
rect 11268 12767 13395 12823
rect 13451 12767 13462 12823
rect 11268 12758 13462 12767
rect 13534 12758 13734 12772
rect 13534 12702 13615 12758
rect 13671 12702 13734 12758
rect 798 12536 2418 12538
rect 798 12492 7646 12536
rect 798 12488 7391 12492
rect 798 12344 852 12488
rect 996 12348 7391 12488
rect 7535 12348 7646 12492
rect 996 12344 7646 12348
rect 798 12300 7646 12344
rect 798 12298 2418 12300
rect 11986 11756 12072 11826
rect 11986 11749 12000 11756
rect 11986 11693 11996 11749
rect 11986 11692 12000 11693
rect 12064 11692 12072 11756
rect 11986 11669 12072 11692
rect 11986 11613 11996 11669
rect 12052 11654 12072 11669
rect 11986 11590 12002 11613
rect 12066 11590 12072 11654
rect 11986 11589 12072 11590
rect 11986 11533 11996 11589
rect 12052 11542 12072 11589
rect 11986 11509 12000 11533
rect 11986 11453 11996 11509
rect 12064 11478 12072 11542
rect 12052 11453 12072 11478
rect 11986 11408 12072 11453
rect 13534 10638 13734 12702
rect 18442 12729 18469 12945
rect 18845 12729 18876 12945
rect 18442 12724 18506 12729
rect 18810 12724 18876 12729
rect 18442 12696 18876 12724
rect 18442 12694 18845 12696
rect 13534 10582 13605 10638
rect 13661 10582 13734 10638
rect 13534 10540 13734 10582
<< via3 >>
rect 8583 38365 8647 38429
rect 5107 33404 5171 33468
rect 5187 33404 5251 33468
rect 5267 33404 5331 33468
rect 7506 33182 7570 33186
rect 7506 33126 7510 33182
rect 7510 33126 7566 33182
rect 7566 33126 7570 33182
rect 7506 33122 7570 33126
rect 7376 33004 7440 33008
rect 7376 32948 7378 33004
rect 7378 32948 7434 33004
rect 7434 32948 7440 33004
rect 7376 32944 7440 32948
rect 9055 31612 9119 31676
rect 23446 33588 23590 33592
rect 23446 33452 23450 33588
rect 23450 33452 23586 33588
rect 23586 33452 23590 33588
rect 23446 33448 23590 33452
rect 16494 31321 16798 31324
rect 849 30730 993 30874
rect 9988 30125 10052 30132
rect 9988 30069 10040 30125
rect 10040 30069 10052 30125
rect 9988 30068 10052 30069
rect 9990 29989 10040 30030
rect 10040 29989 10054 30030
rect 9990 29966 10054 29989
rect 9988 29909 10040 29918
rect 10040 29909 10052 29918
rect 9988 29885 10052 29909
rect 9988 29854 10040 29885
rect 10040 29854 10052 29885
rect 16494 31105 16798 31321
rect 16494 31100 16798 31105
rect 10602 19902 10666 19966
rect 25732 19116 25796 19120
rect 25732 19060 25736 19116
rect 25736 19060 25792 19116
rect 25792 19060 25796 19116
rect 25732 19056 25796 19060
rect 10602 15278 10666 15282
rect 10602 15222 10606 15278
rect 10606 15222 10662 15278
rect 10662 15222 10666 15278
rect 10602 15218 10666 15222
rect 9517 14806 9581 14810
rect 9517 14750 9521 14806
rect 9521 14750 9577 14806
rect 9577 14750 9581 14806
rect 9517 14746 9581 14750
rect 9388 14628 9452 14632
rect 9388 14572 9390 14628
rect 9390 14572 9446 14628
rect 9446 14572 9452 14628
rect 9388 14568 9452 14572
rect 10882 13732 10946 13796
rect 25458 15212 25602 15216
rect 25458 15076 25462 15212
rect 25462 15076 25598 15212
rect 25598 15076 25602 15212
rect 25458 15072 25602 15076
rect 18506 12945 18810 12948
rect 7391 12489 7535 12492
rect 852 12344 996 12488
rect 7391 12353 7396 12489
rect 7396 12353 7532 12489
rect 7532 12353 7535 12489
rect 7391 12348 7535 12353
rect 12000 11749 12064 11756
rect 12000 11693 12052 11749
rect 12052 11693 12064 11749
rect 12000 11692 12064 11693
rect 12002 11613 12052 11654
rect 12052 11613 12066 11654
rect 12002 11590 12066 11613
rect 12000 11533 12052 11542
rect 12052 11533 12064 11542
rect 12000 11509 12064 11533
rect 12000 11478 12052 11509
rect 12052 11478 12064 11509
rect 18506 12729 18810 12945
rect 18506 12724 18810 12729
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 200 1000 440 44152
rect 800 30874 1040 44152
rect 800 30730 849 30874
rect 993 30730 1040 30874
rect 800 12488 1040 30730
rect 800 12344 852 12488
rect 996 12344 1040 12488
rect 800 1000 1040 12344
rect 1600 33478 1840 44152
rect 11341 43905 11441 44005
rect 11341 43805 11541 43905
rect 11721 43897 11835 44009
rect 11615 43805 11835 43897
rect 11341 43705 11835 43805
rect 11341 43305 11441 43705
rect 11541 43697 11835 43705
rect 11541 43605 11641 43697
rect 11721 43309 11835 43697
rect 11913 43927 12401 44013
rect 11913 43725 12027 43927
rect 12287 43725 12401 43927
rect 11913 43639 12401 43725
rect 11913 43313 12027 43639
rect 12287 43313 12401 43639
rect 12611 43905 12711 44005
rect 12611 43805 12811 43905
rect 12991 43897 13105 44009
rect 12885 43805 13105 43897
rect 12611 43705 13105 43805
rect 12611 43305 12711 43705
rect 12811 43697 13105 43705
rect 12811 43605 12911 43697
rect 12991 43309 13105 43697
rect 13171 43927 13615 44013
rect 13171 43711 13285 43927
rect 13735 43905 14135 44005
rect 13171 43625 13613 43711
rect 13171 43399 13285 43625
rect 13735 43405 13835 43905
rect 14035 43805 14235 43905
rect 14135 43505 14235 43805
rect 14035 43405 14235 43505
rect 14329 43697 14429 43997
rect 14629 43697 14729 43997
rect 14329 43597 14729 43697
rect 13169 43313 13611 43399
rect 13735 43305 14135 43405
rect 14329 43297 14429 43597
rect 14629 43297 14729 43597
rect 14829 43913 15317 43999
rect 14829 43711 14943 43913
rect 15203 43711 15317 43913
rect 14829 43625 15317 43711
rect 14829 43299 14943 43625
rect 15203 43299 15317 43625
rect 9321 42083 9521 42883
rect 10221 42683 10921 42883
rect 10221 42483 10421 42683
rect 10721 42483 10921 42683
rect 10221 42283 10921 42483
rect 11121 42683 11821 42883
rect 12021 42683 12721 42883
rect 9321 41883 10021 42083
rect 10221 41883 10421 42283
rect 11121 42083 11321 42683
rect 12021 42483 12221 42683
rect 12521 42483 12721 42683
rect 12021 42283 12721 42483
rect 12921 42683 13621 42883
rect 12921 42483 13121 42683
rect 12921 42283 13621 42483
rect 14021 42283 14521 42483
rect 11121 41883 11821 42083
rect 12021 41883 12221 42283
rect 12521 41883 12721 42283
rect 13421 42083 13621 42283
rect 12921 41883 13621 42083
rect 14721 41883 14921 42883
rect 15121 41883 15321 42883
rect 15521 42683 16321 42883
rect 16521 42683 17321 42883
rect 17521 42783 17721 42883
rect 15821 41883 16021 42683
rect 16521 42083 16721 42683
rect 17521 42583 17921 42783
rect 16921 42283 17321 42483
rect 17121 42083 17321 42283
rect 16521 41883 17321 42083
rect 17521 41883 17721 42583
rect 17821 42483 18021 42583
rect 17921 42383 18121 42483
rect 18021 42283 18221 42383
rect 18321 42283 18521 42883
rect 18121 42183 18521 42283
rect 18221 42083 18521 42183
rect 18321 41883 18521 42083
rect 8546 40750 8646 40850
rect 8546 40650 8746 40750
rect 8546 40550 8846 40650
rect 8546 40150 8646 40550
rect 8746 40450 8946 40550
rect 9046 40450 9146 40850
rect 8846 40350 9146 40450
rect 8946 40250 9146 40350
rect 9046 40150 9146 40250
rect 9246 40150 9346 40850
rect 9446 40750 9946 40850
rect 9646 40150 9746 40750
rect 10046 40550 10146 40850
rect 10446 40550 10546 40850
rect 10046 40450 10546 40550
rect 10046 40150 10146 40450
rect 10446 40150 10546 40450
rect 10646 40150 10746 40850
rect 10846 40750 10946 40850
rect 10846 40650 11046 40750
rect 10846 40550 11146 40650
rect 10846 40150 10946 40550
rect 11046 40450 11246 40550
rect 11346 40450 11446 40850
rect 11146 40350 11446 40450
rect 11246 40250 11446 40350
rect 11346 40150 11446 40250
rect 11646 40750 12046 40850
rect 11646 40550 11746 40750
rect 11946 40550 12046 40750
rect 11646 40450 12046 40550
rect 12546 40550 12646 40850
rect 12946 40750 13046 40850
rect 12846 40650 13046 40750
rect 13146 40750 13546 40850
rect 12746 40550 12946 40650
rect 13146 40550 13246 40750
rect 13446 40550 13546 40750
rect 12546 40450 12846 40550
rect 13146 40450 13546 40550
rect 11646 40150 11746 40450
rect 12546 40150 12646 40450
rect 12746 40350 12946 40450
rect 12846 40250 13046 40350
rect 12946 40150 13046 40250
rect 13146 40150 13246 40450
rect 13446 40150 13546 40450
rect 13646 40750 14046 40850
rect 14146 40750 14646 40850
rect 13646 40550 13746 40750
rect 13946 40550 14046 40750
rect 13646 40450 14046 40550
rect 13646 40150 13746 40450
rect 13846 40350 13946 40450
rect 13846 40250 14046 40350
rect 13946 40150 14046 40250
rect 14346 40150 14446 40750
rect 14746 40150 14846 40850
rect 14946 40550 15046 40850
rect 15346 40750 15446 40850
rect 15246 40650 15446 40750
rect 15546 40750 15946 40850
rect 15146 40550 15346 40650
rect 15546 40550 15646 40750
rect 15846 40550 15946 40750
rect 14946 40450 15246 40550
rect 15546 40450 15946 40550
rect 16046 40550 16146 40850
rect 16346 40550 16446 40850
rect 16046 40450 16446 40550
rect 16946 40750 17146 40850
rect 17446 40750 17646 40850
rect 16946 40650 17246 40750
rect 17346 40650 17646 40750
rect 14946 40150 15046 40450
rect 15146 40350 15346 40450
rect 15246 40250 15446 40350
rect 15346 40150 15446 40250
rect 15546 40150 15646 40450
rect 15846 40150 15946 40450
rect 16196 40150 16296 40450
rect 16946 40150 17046 40650
rect 17146 40550 17646 40650
rect 17246 40450 17346 40550
rect 17546 40150 17646 40550
rect 17746 40750 18146 40850
rect 17746 40550 17846 40750
rect 18046 40550 18146 40750
rect 17746 40450 18146 40550
rect 17746 40150 17846 40450
rect 18046 40150 18146 40450
rect 18246 40750 18646 40850
rect 18246 40250 18346 40750
rect 18546 40650 18746 40750
rect 18646 40350 18746 40650
rect 18546 40250 18746 40350
rect 18846 40550 18946 40850
rect 19146 40550 19246 40850
rect 18846 40450 19246 40550
rect 18246 40150 18646 40250
rect 18846 40150 18946 40450
rect 19146 40150 19246 40450
rect 19346 40750 19746 40850
rect 19346 40550 19446 40750
rect 19646 40550 19746 40750
rect 19346 40450 19746 40550
rect 19346 40150 19446 40450
rect 19646 40150 19746 40450
rect 19846 40450 19946 40850
rect 20346 40450 20446 40850
rect 19846 40350 20046 40450
rect 20246 40350 20446 40450
rect 20646 40750 21146 40850
rect 20646 40550 20746 40750
rect 20946 40550 21146 40750
rect 20646 40450 21146 40550
rect 19946 40250 20346 40350
rect 20046 40150 20246 40250
rect 20646 40150 20746 40450
rect 22878 38462 22938 45152
rect 8566 38429 22938 38462
rect 8566 38365 8583 38429
rect 8647 38365 22938 38429
rect 8566 38340 22938 38365
rect 8566 38330 22936 38340
rect 8566 38328 9094 38330
rect 23430 37872 23490 45152
rect 7478 37758 23490 37872
rect 1600 33468 5386 33478
rect 1600 33404 5107 33468
rect 5171 33404 5187 33468
rect 5251 33404 5267 33468
rect 5331 33404 5386 33468
rect 1600 33394 5386 33404
rect 1600 1000 1840 33394
rect 7480 33186 7596 37758
rect 7480 33122 7506 33186
rect 7570 33122 7596 33186
rect 7480 33098 7596 33122
rect 23356 33592 23788 33658
rect 23356 33448 23446 33592
rect 23590 33448 23788 33592
rect 7356 33036 21286 33038
rect 23356 33036 23788 33448
rect 7356 33034 23788 33036
rect 7356 33008 23782 33034
rect 7356 32944 7376 33008
rect 7440 32944 23782 33008
rect 7356 32922 23782 32944
rect 7328 12492 7646 12536
rect 7328 12348 7391 12492
rect 7535 12348 7646 12492
rect 7328 12300 7646 12348
rect 7914 984 8094 32922
rect 9008 31682 9100 31684
rect 9008 31676 9166 31682
rect 9008 31612 9055 31676
rect 9119 31612 9166 31676
rect 9008 1600 9166 31612
rect 16434 31384 18694 31388
rect 16326 31324 18694 31384
rect 16326 31100 16494 31324
rect 16798 31100 18694 31324
rect 16326 31050 18694 31100
rect 16328 30818 16430 31050
rect 18588 30804 18694 31050
rect 9984 30132 16002 30202
rect 9984 30068 9988 30132
rect 10052 30068 16002 30132
rect 9984 30030 16002 30068
rect 9984 29966 9990 30030
rect 10054 29966 16002 30030
rect 9984 29918 16002 29966
rect 9984 29854 9988 29918
rect 10052 29854 16002 29918
rect 9984 29784 16002 29854
rect 15220 22860 15326 23096
rect 17482 22860 17588 23140
rect 15220 22766 17588 22860
rect 10582 19984 10686 19988
rect 23982 19984 24042 45152
rect 10582 19966 24042 19984
rect 10582 19902 10602 19966
rect 10666 19902 24042 19966
rect 10582 19884 24042 19902
rect 24534 19626 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 9496 19522 24594 19626
rect 9496 18204 9596 19522
rect 27234 19136 27414 19380
rect 25714 19120 27414 19136
rect 25714 19056 25732 19120
rect 25796 19056 27414 19120
rect 25714 19038 27414 19056
rect 9496 14810 9602 18204
rect 10584 15282 10682 15312
rect 10584 15218 10602 15282
rect 10666 15218 10682 15282
rect 10584 15202 10682 15218
rect 25368 15216 25800 15282
rect 9496 14746 9517 14810
rect 9581 14746 9602 14810
rect 9496 14726 9602 14746
rect 25368 15072 25458 15216
rect 25602 15072 25800 15216
rect 9368 14660 23298 14662
rect 25368 14660 25800 15072
rect 9368 14658 25800 14660
rect 9368 14632 25794 14658
rect 9368 14568 9388 14632
rect 9452 14568 25794 14632
rect 9368 14546 25794 14568
rect 10862 13796 10966 13824
rect 10862 13732 10882 13796
rect 10946 13732 10966 13796
rect 10862 2054 10966 13732
rect 19506 13012 19686 14546
rect 18446 13008 20706 13012
rect 18338 12948 20706 13008
rect 18338 12724 18506 12948
rect 18810 12724 20706 12948
rect 18338 12674 20706 12724
rect 18340 12442 18442 12674
rect 11996 11756 18014 11826
rect 11996 11692 12000 11756
rect 12064 11692 18014 11756
rect 11996 11654 18014 11692
rect 11996 11590 12002 11654
rect 12066 11590 18014 11654
rect 11996 11542 18014 11590
rect 11996 11478 12000 11542
rect 12064 11478 18014 11542
rect 11996 11408 18014 11478
rect 19506 4764 19686 12674
rect 20600 12428 20706 12674
rect 17232 4484 17338 4720
rect 19494 4484 19686 4764
rect 17232 4390 19686 4484
rect 10860 1830 19686 2054
rect 10860 1828 11214 1830
rect 15568 1600 15822 1602
rect 9008 1598 11220 1600
rect 12160 1598 15822 1600
rect 9008 1420 15822 1598
rect 9190 984 11958 986
rect 7912 824 11958 984
rect 9190 820 11958 824
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 820
rect 15642 0 15822 1420
rect 19506 0 19686 1830
rect 23370 0 23550 14546
rect 27234 0 27414 19038
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_0
timestamp 1748330293
transform 1 0 12726 0 1 12270
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_1
timestamp 1748330293
transform 1 0 12014 0 1 12116
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_2
timestamp 1748330293
transform 1 0 12726 0 1 13448
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_3
timestamp 1748330293
transform 1 0 12014 0 1 13606
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_4
timestamp 1748330293
transform 1 0 10002 0 1 30492
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_5
timestamp 1748330293
transform 1 0 10714 0 1 30646
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_6
timestamp 1748330293
transform 1 0 10714 0 1 31824
box -23 -33 23 33
use L1M1_C_CDNS_741011383740  L1M1_C_CDNS_741011383740_7
timestamp 1748330293
transform 1 0 10002 0 1 31982
box -23 -33 23 33
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_0
timestamp 1748330293
transform 1 0 11658 0 1 12515
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_1
timestamp 1748330293
transform 1 0 12370 0 1 12515
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_2
timestamp 1748330293
transform 1 0 13082 0 1 12515
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_3
timestamp 1748330293
transform 1 0 11658 0 1 13207
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_4
timestamp 1748330293
transform 1 0 12370 0 1 13207
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_5
timestamp 1748330293
transform 1 0 13082 0 1 13207
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_6
timestamp 1748330293
transform 1 0 12262 0 1 17623
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_7
timestamp 1748330293
transform 1 0 14336 0 1 17623
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_8
timestamp 1748330293
transform 1 0 14760 0 1 15426
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_9
timestamp 1748330293
transform 1 0 15647 0 1 18099
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_10
timestamp 1748330293
transform 1 0 13025 0 1 18099
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_11
timestamp 1748330293
transform 1 0 9646 0 1 31583
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_12
timestamp 1748330293
transform 1 0 9646 0 1 30891
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_13
timestamp 1748330293
transform 1 0 10358 0 1 31583
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_14
timestamp 1748330293
transform 1 0 10358 0 1 30891
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_15
timestamp 1748330293
transform 1 0 11070 0 1 31583
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_16
timestamp 1748330293
transform 1 0 11070 0 1 30891
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_17
timestamp 1748330293
transform 1 0 12748 0 1 33802
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_18
timestamp 1748330293
transform 1 0 10250 0 1 35999
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_19
timestamp 1748330293
transform 1 0 12324 0 1 35999
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_20
timestamp 1748330293
transform 1 0 13635 0 1 36475
box -23 -105 23 105
use L1M1_C_CDNS_741011383742  L1M1_C_CDNS_741011383742_21
timestamp 1748330293
transform 1 0 11013 0 1 36475
box -23 -105 23 105
use L1M1_C_CDNS_741011383743  L1M1_C_CDNS_741011383743_0
timestamp 1748330293
transform 1 0 16410 0 1 17623
box -23 -101 23 101
use L1M1_C_CDNS_741011383743  L1M1_C_CDNS_741011383743_1
timestamp 1748330293
transform 1 0 14248 0 1 15426
box -23 -101 23 101
use L1M1_C_CDNS_741011383743  L1M1_C_CDNS_741011383743_2
timestamp 1748330293
transform 1 0 12236 0 1 33802
box -23 -101 23 101
use L1M1_C_CDNS_741011383743  L1M1_C_CDNS_741011383743_3
timestamp 1748330293
transform 1 0 14398 0 1 35999
box -23 -101 23 101
use L1M1_C_CDNS_7410113837410  L1M1_C_CDNS_7410113837410_0
timestamp 1748330293
transform 1 0 14591 0 -1 13946
box -23 -37 23 37
use L1M1_C_CDNS_7410113837410  L1M1_C_CDNS_7410113837410_1
timestamp 1748330293
transform 1 0 20460 0 1 17616
box -23 -37 23 37
use L1M1_C_CDNS_7410113837410  L1M1_C_CDNS_7410113837410_2
timestamp 1748330293
transform 1 0 12579 0 -1 32322
box -23 -37 23 37
use L1M1_C_CDNS_7410113837410  L1M1_C_CDNS_7410113837410_3
timestamp 1748330293
transform 1 0 18448 0 1 35992
box -23 -37 23 37
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_0
timestamp 1748330293
transform 1 0 17131 0 -1 13946
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_1
timestamp 1748330293
transform 1 0 25708 0 1 17616
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_2
timestamp 1748330293
transform 1 0 23084 0 1 17616
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_3
timestamp 1748330293
transform 1 0 20070 0 1 17614
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_4
timestamp 1748330293
transform 1 0 15119 0 -1 32322
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_5
timestamp 1748330293
transform 1 0 18058 0 1 35990
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_6
timestamp 1748330293
transform 1 0 21072 0 1 35992
box -32 -26 32 26
use L1M1_C_CDNS_7410113837414  L1M1_C_CDNS_7410113837414_7
timestamp 1748330293
transform 1 0 23696 0 1 35992
box -32 -26 32 26
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_0
timestamp 1748330293
transform 1 0 11883 0 1 31216
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_1
timestamp 1748330293
transform 1 0 16090 0 1 35990
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_2
timestamp 1748330293
transform 1 0 21116 0 1 17615
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_3
timestamp 1748330293
transform 1 0 18102 0 1 17614
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_4
timestamp 1748330293
transform 1 0 19414 0 1 17614
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_5
timestamp 1748330293
transform 1 0 13895 0 1 12840
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_6
timestamp 1748330293
transform 1 0 17402 0 1 35990
box -29 -23 29 23
use L1M1_C_CDNS_7410113837415  L1M1_C_CDNS_7410113837415_7
timestamp 1748330293
transform 1 0 19104 0 1 35991
box -29 -23 29 23
use L1M1_C_CDNS_7410113837416  L1M1_C_CDNS_7410113837416_0
timestamp 1748330293
transform 1 0 22428 0 1 17615
box -23 -29 23 29
use L1M1_C_CDNS_7410113837416  L1M1_C_CDNS_7410113837416_1
timestamp 1748330293
transform 1 0 20416 0 1 35991
box -23 -29 23 29
use L1M1_C_CDNS_7410113837417  L1M1_C_CDNS_7410113837417_0
timestamp 1748330293
transform 1 0 17446 0 1 17614
box -37 -23 37 23
use L1M1_C_CDNS_7410113837417  L1M1_C_CDNS_7410113837417_1
timestamp 1748330293
transform 1 0 15434 0 1 35990
box -37 -23 37 23
use L1M1_C_CDNS_7410113837422  L1M1_C_CDNS_7410113837422_0
timestamp 1748330293
transform 1 0 12678 0 1 15252
box -26 -128 26 128
use L1M1_C_CDNS_7410113837422  L1M1_C_CDNS_7410113837422_1
timestamp 1748330293
transform 1 0 10666 0 1 33628
box -26 -128 26 128
use L1M1_C_CDNS_7410113837423  L1M1_C_CDNS_7410113837423_0
timestamp 1748330293
transform 1 0 15904 0 1 15471
box -23 -245 23 245
use L1M1_C_CDNS_7410113837423  L1M1_C_CDNS_7410113837423_1
timestamp 1748330293
transform 1 0 13892 0 1 33847
box -23 -245 23 245
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_0
timestamp 1748330293
transform 1 0 11606 0 1 16913
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_1
timestamp 1748330293
transform 1 0 12370 0 1 16604
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_2
timestamp 1748330293
transform 1 0 17025 0 1 14184
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_3
timestamp 1748330293
transform 1 0 16302 0 1 16604
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_4
timestamp 1748330293
transform 1 0 9594 0 1 35289
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_5
timestamp 1748330293
transform 1 0 10358 0 1 34980
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_6
timestamp 1748330293
transform 1 0 15013 0 1 32560
box -26 -32 26 32
use L1M1_C_CDNS_7410113837436  L1M1_C_CDNS_7410113837436_7
timestamp 1748330293
transform 1 0 14290 0 1 34980
box -26 -32 26 32
use L1M1_C_CDNS_7410113837450  L1M1_C_CDNS_7410113837450_0
timestamp 1748330293
transform 1 0 21421 0 1 15717
box -23 -100 23 100
use L1M1_C_CDNS_7410113837450  L1M1_C_CDNS_7410113837450_1
timestamp 1748330293
transform 1 0 19409 0 1 34093
box -23 -100 23 100
use L1M1_C_CDNS_7410113837456  L1M1_C_CDNS_7410113837456_0
timestamp 1748330293
transform 1 0 20070 0 1 16293
box -23 -65 23 65
use L1M1_C_CDNS_7410113837456  L1M1_C_CDNS_7410113837456_1
timestamp 1748330293
transform 1 0 18058 0 1 34669
box -23 -65 23 65
use L1M1_C_CDNS_7410113837457  L1M1_C_CDNS_7410113837457_0
timestamp 1748330293
transform 1 0 25708 0 1 16585
box -23 -353 23 353
use L1M1_C_CDNS_7410113837457  L1M1_C_CDNS_7410113837457_1
timestamp 1748330293
transform 1 0 23696 0 1 34961
box -23 -353 23 353
use L1M1_C_CDNS_7410113837460  L1M1_C_CDNS_7410113837460_0
timestamp 1748330293
transform 1 0 13639 0 1 12754
box -68 -23 68 23
use L1M1_C_CDNS_7410113837460  L1M1_C_CDNS_7410113837460_1
timestamp 1748330293
transform 1 0 11627 0 1 31130
box -68 -23 68 23
use L1M1_C_CDNS_7410113837463  L1M1_C_CDNS_7410113837463_0
timestamp 1748330293
transform 1 0 17083 0 1 16913
box -43 -32 9 32
use L1M1_C_CDNS_7410113837463  L1M1_C_CDNS_7410113837463_1
timestamp 1748330293
transform 1 0 15071 0 1 35289
box -43 -32 9 32
use L1M1_C_CDNS_7410113837465  L1M1_C_CDNS_7410113837465_0
timestamp 1748330293
transform 1 0 9204 0 1 14581
box -37 -29 37 17
use L1M1_C_CDNS_7410113837465  L1M1_C_CDNS_7410113837465_1
timestamp 1748330293
transform 1 0 7192 0 1 32957
box -37 -29 37 17
use L1M1_C_CDNS_7410113837467  L1M1_C_CDNS_7410113837467_0
timestamp 1748330293
transform 1 0 9921 0 1 15144
box -29 -27 29 27
use L1M1_C_CDNS_7410113837467  L1M1_C_CDNS_7410113837467_1
timestamp 1748330293
transform 1 0 7909 0 1 33520
box -29 -27 29 27
use L1M1_C_CDNS_7410113837468  L1M1_C_CDNS_7410113837468_0
timestamp 1748330293
transform 1 0 11379 0 1 14416
box -29 -27 29 27
use L1M1_C_CDNS_7410113837468  L1M1_C_CDNS_7410113837468_1
timestamp 1748330293
transform 1 0 9367 0 1 32792
box -29 -27 29 27
use L1M1_C_CDNS_7410113837471  L1M1_C_CDNS_7410113837471_0
timestamp 1748330293
transform 1 0 9793 0 1 14611
box -55 -23 55 23
use L1M1_C_CDNS_7410113837471  L1M1_C_CDNS_7410113837471_1
timestamp 1748330293
transform 1 0 7781 0 1 32987
box -55 -23 55 23
use L1M1_C_CDNS_7410113837472  L1M1_C_CDNS_7410113837472_0
timestamp 1748330293
transform 1 0 9759 0 1 14986
box -55 -15 55 31
use L1M1_C_CDNS_7410113837472  L1M1_C_CDNS_7410113837472_1
timestamp 1748330293
transform 1 0 7747 0 1 33362
box -55 -15 55 31
use L1M1_C_CDNS_7410113837473  L1M1_C_CDNS_7410113837473_0
timestamp 1748330293
transform 1 0 9513 0 1 13387
box -23 -51 23 51
use L1M1_C_CDNS_7410113837473  L1M1_C_CDNS_7410113837473_1
timestamp 1748330293
transform 1 0 7501 0 1 31763
box -23 -51 23 51
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_0
timestamp 1748330293
transform 1 0 12734 0 1 12769
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_1
timestamp 1748330293
transform 1 0 12013 0 1 12953
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_2
timestamp 1748330293
transform 1 0 11713 0 1 12953
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_3
timestamp 1748330293
transform 1 0 13027 0 1 12953
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_4
timestamp 1748330293
transform 1 0 11713 0 1 11035
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_5
timestamp 1748330293
transform 1 0 9701 0 1 29411
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_6
timestamp 1748330293
transform 1 0 9701 0 1 31329
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_7
timestamp 1748330293
transform 1 0 10001 0 1 31329
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_8
timestamp 1748330293
transform 1 0 11015 0 1 31329
box -32 -32 32 32
use M1M2_C_CDNS_741011383741  M1M2_C_CDNS_741011383741_9
timestamp 1748330293
transform 1 0 10722 0 1 31145
box -32 -32 32 32
use M1M2_C_CDNS_741011383744  M1M2_C_CDNS_741011383744_0
timestamp 1748330293
transform 1 0 12913 0 1 16173
box -64 -27 64 27
use M1M2_C_CDNS_741011383744  M1M2_C_CDNS_741011383744_1
timestamp 1748330293
transform 1 0 12785 0 1 16173
box -64 -27 64 27
use M1M2_C_CDNS_741011383744  M1M2_C_CDNS_741011383744_2
timestamp 1748330293
transform 1 0 10773 0 1 34549
box -64 -27 64 27
use M1M2_C_CDNS_741011383744  M1M2_C_CDNS_741011383744_3
timestamp 1748330293
transform 1 0 10901 0 1 34549
box -64 -27 64 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_0
timestamp 1748330293
transform 1 0 15834 0 1 16173
box -128 -27 128 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_1
timestamp 1748330293
transform -1 0 19591 0 1 16173
box -128 -27 128 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_2
timestamp 1748330293
transform -1 0 17928 0 1 16173
box -128 -27 128 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_3
timestamp 1748330293
transform 1 0 13822 0 1 34549
box -128 -27 128 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_4
timestamp 1748330293
transform -1 0 15916 0 1 34549
box -128 -27 128 27
use M1M2_C_CDNS_741011383745  M1M2_C_CDNS_741011383745_5
timestamp 1748330293
transform -1 0 17579 0 1 34549
box -128 -27 128 27
use M1M2_C_CDNS_741011383746  M1M2_C_CDNS_741011383746_0
timestamp 1748330293
transform -1 0 22643 0 1 16173
box -160 -27 160 27
use M1M2_C_CDNS_741011383746  M1M2_C_CDNS_741011383746_1
timestamp 1748330293
transform -1 0 20918 0 1 16173
box -160 -27 160 27
use M1M2_C_CDNS_741011383746  M1M2_C_CDNS_741011383746_2
timestamp 1748330293
transform -1 0 18906 0 1 34549
box -160 -27 160 27
use M1M2_C_CDNS_741011383746  M1M2_C_CDNS_741011383746_3
timestamp 1748330293
transform -1 0 20631 0 1 34549
box -160 -27 160 27
use M1M2_C_CDNS_7410113837412  M1M2_C_CDNS_7410113837412_0
timestamp 1748330293
transform 1 0 14591 0 -1 13946
box -32 -37 32 37
use M1M2_C_CDNS_7410113837412  M1M2_C_CDNS_7410113837412_1
timestamp 1748330293
transform 1 0 20460 0 1 17616
box -32 -37 32 37
use M1M2_C_CDNS_7410113837412  M1M2_C_CDNS_7410113837412_2
timestamp 1748330293
transform 1 0 12579 0 -1 32322
box -32 -37 32 37
use M1M2_C_CDNS_7410113837412  M1M2_C_CDNS_7410113837412_3
timestamp 1748330293
transform 1 0 18448 0 1 35992
box -32 -37 32 37
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_0
timestamp 1748330293
transform 1 0 17131 0 -1 13946
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_1
timestamp 1748330293
transform 1 0 25708 0 1 17616
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_2
timestamp 1748330293
transform 1 0 23084 0 1 17616
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_3
timestamp 1748330293
transform 1 0 20070 0 1 17614
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_4
timestamp 1748330293
transform 1 0 15119 0 -1 32322
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_5
timestamp 1748330293
transform 1 0 18058 0 1 35990
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_6
timestamp 1748330293
transform 1 0 21072 0 1 35992
box -32 -26 32 26
use M1M2_C_CDNS_7410113837413  M1M2_C_CDNS_7410113837413_7
timestamp 1748330293
transform 1 0 23696 0 1 35992
box -32 -26 32 26
use M1M2_C_CDNS_7410113837418  M1M2_C_CDNS_7410113837418_0
timestamp 1748330293
transform 1 0 12806 0 1 15057
box -96 -26 96 26
use M1M2_C_CDNS_7410113837418  M1M2_C_CDNS_7410113837418_1
timestamp 1748330293
transform 1 0 10794 0 1 33433
box -96 -26 96 26
use M1M2_C_CDNS_7410113837419  M1M2_C_CDNS_7410113837419_0
timestamp 1748330293
transform 1 0 17446 0 1 17614
box -37 -26 37 26
use M1M2_C_CDNS_7410113837419  M1M2_C_CDNS_7410113837419_1
timestamp 1748330293
transform 1 0 15434 0 1 35990
box -37 -26 37 26
use M1M2_C_CDNS_7410113837420  M1M2_C_CDNS_7410113837420_0
timestamp 1748330293
transform 1 0 11548 0 1 14393
box -26 -32 26 32
use M1M2_C_CDNS_7410113837420  M1M2_C_CDNS_7410113837420_1
timestamp 1748330293
transform 1 0 13196 0 1 14002
box -26 -32 26 32
use M1M2_C_CDNS_7410113837420  M1M2_C_CDNS_7410113837420_2
timestamp 1748330293
transform 1 0 9536 0 1 32769
box -26 -32 26 32
use M1M2_C_CDNS_7410113837420  M1M2_C_CDNS_7410113837420_3
timestamp 1748330293
transform 1 0 11184 0 1 32378
box -26 -32 26 32
use M1M2_C_CDNS_7410113837421  M1M2_C_CDNS_7410113837421_0
timestamp 1748330293
transform 1 0 12678 0 1 15252
box -26 -128 26 128
use M1M2_C_CDNS_7410113837421  M1M2_C_CDNS_7410113837421_1
timestamp 1748330293
transform 1 0 10666 0 1 33628
box -26 -128 26 128
use M1M2_C_CDNS_7410113837424  M1M2_C_CDNS_7410113837424_0
timestamp 1748330293
transform 1 0 15904 0 1 15471
box -26 -256 26 256
use M1M2_C_CDNS_7410113837424  M1M2_C_CDNS_7410113837424_1
timestamp 1748330293
transform 1 0 13892 0 1 33847
box -26 -256 26 256
use M1M2_C_CDNS_7410113837425  M1M2_C_CDNS_7410113837425_0
timestamp 1748330293
transform 1 0 16147 0 1 14537
box -160 -26 160 26
use M1M2_C_CDNS_7410113837425  M1M2_C_CDNS_7410113837425_1
timestamp 1748330293
transform 1 0 14135 0 1 32913
box -160 -26 160 26
use M1M2_C_CDNS_7410113837426  M1M2_C_CDNS_7410113837426_0
timestamp 1748330293
transform 1 0 15572 0 1 14537
box -192 -26 192 26
use M1M2_C_CDNS_7410113837427  M1M2_C_CDNS_7410113837427_0
timestamp 1748330293
transform 1 0 14591 0 1 15426
box -32 -101 32 101
use M1M2_C_CDNS_7410113837427  M1M2_C_CDNS_7410113837427_1
timestamp 1748330293
transform 1 0 12579 0 1 33802
box -32 -101 32 101
use M1M2_C_CDNS_7410113837429  M1M2_C_CDNS_7410113837429_0
timestamp 1748330293
transform 1 0 14469 0 1 15660
box -101 -90 101 90
use M1M2_C_CDNS_7410113837429  M1M2_C_CDNS_7410113837429_1
timestamp 1748330293
transform 1 0 14469 0 1 15995
box -101 -90 101 90
use M1M2_C_CDNS_7410113837429  M1M2_C_CDNS_7410113837429_2
timestamp 1748330293
transform 1 0 12457 0 1 34036
box -101 -90 101 90
use M1M2_C_CDNS_7410113837429  M1M2_C_CDNS_7410113837429_3
timestamp 1748330293
transform 1 0 12457 0 1 34371
box -101 -90 101 90
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_0
timestamp 1748330293
transform 1 0 12370 0 1 16603
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_1
timestamp 1748330293
transform 1 0 11606 0 1 16913
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_2
timestamp 1748330293
transform 1 0 17025 0 1 14184
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_3
timestamp 1748330293
transform 1 0 21378 0 1 15915
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_4
timestamp 1748330293
transform 1 0 16304 0 1 16607
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_5
timestamp 1748330293
transform 1 0 9594 0 1 35289
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_6
timestamp 1748330293
transform 1 0 10358 0 1 34979
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_7
timestamp 1748330293
transform 1 0 15013 0 1 32560
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_8
timestamp 1748330293
transform 1 0 14292 0 1 34983
box -28 -37 28 37
use M1M2_C_CDNS_7410113837435  M1M2_C_CDNS_7410113837435_9
timestamp 1748330293
transform 1 0 19366 0 1 34291
box -28 -37 28 37
use M1M2_C_CDNS_7410113837446  M1M2_C_CDNS_7410113837446_0
timestamp 1748330293
transform 1 0 21773 0 1 16065
box -32 -32 32 32
use M1M2_C_CDNS_7410113837446  M1M2_C_CDNS_7410113837446_1
timestamp 1748330293
transform 1 0 18760 0 1 16065
box -32 -32 32 32
use M1M2_C_CDNS_7410113837446  M1M2_C_CDNS_7410113837446_2
timestamp 1748330293
transform 1 0 16748 0 1 34441
box -32 -32 32 32
use M1M2_C_CDNS_7410113837446  M1M2_C_CDNS_7410113837446_3
timestamp 1748330293
transform 1 0 19761 0 1 34441
box -32 -32 32 32
use M1M2_C_CDNS_7410113837447  M1M2_C_CDNS_7410113837447_0
timestamp 1748330293
transform 1 0 14115 0 1 14973
box -32 -32 32 32
use M1M2_C_CDNS_7410113837447  M1M2_C_CDNS_7410113837447_1
timestamp 1748330293
transform 1 0 12103 0 1 33349
box -32 -32 32 32
use M1M2_C_CDNS_7410113837454  M1M2_C_CDNS_7410113837454_0
timestamp 1748330293
transform 1 0 25708 0 1 16585
box -26 -353 26 353
use M1M2_C_CDNS_7410113837454  M1M2_C_CDNS_7410113837454_1
timestamp 1748330293
transform 1 0 23696 0 1 34961
box -26 -353 26 353
use M1M2_C_CDNS_7410113837458  M1M2_C_CDNS_7410113837458_0
timestamp 1748330293
transform 1 0 20070 0 1 16293
box -26 -65 26 65
use M1M2_C_CDNS_7410113837458  M1M2_C_CDNS_7410113837458_1
timestamp 1748330293
transform 1 0 18058 0 1 34669
box -26 -65 26 65
use M1M2_C_CDNS_7410113837462  M1M2_C_CDNS_7410113837462_0
timestamp 1748330293
transform 1 0 17083 0 1 16913
box -45 -37 11 37
use M1M2_C_CDNS_7410113837462  M1M2_C_CDNS_7410113837462_1
timestamp 1748330293
transform 1 0 15071 0 1 35289
box -45 -37 11 37
use M1M2_C_CDNS_7410113837466  M1M2_C_CDNS_7410113837466_0
timestamp 1748330293
transform 1 0 9204 0 1 14581
box -50 -32 50 20
use M1M2_C_CDNS_7410113837466  M1M2_C_CDNS_7410113837466_1
timestamp 1748330293
transform 1 0 7192 0 1 32957
box -50 -32 50 20
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_0
timestamp 1748330293
transform 1 0 11713 0 1 14741
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_1
timestamp 1748330293
transform 1 0 11606 0 1 16913
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_2
timestamp 1748330293
transform 1 0 13027 0 1 14743
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_3
timestamp 1748330293
transform 1 0 12369 0 1 16603
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_4
timestamp 1748330293
transform 1 0 16309 0 1 16599
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_5
timestamp 1748330293
transform 1 0 17025 0 1 14184
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_6
timestamp 1748330293
transform 1 0 21378 0 1 15915
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_7
timestamp 1748330293
transform 1 0 9701 0 1 33117
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_8
timestamp 1748330293
transform 1 0 9594 0 1 35289
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_9
timestamp 1748330293
transform 1 0 11015 0 1 33119
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_10
timestamp 1748330293
transform 1 0 10357 0 1 34979
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_11
timestamp 1748330293
transform 1 0 15013 0 1 32560
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_12
timestamp 1748330293
transform 1 0 14297 0 1 34975
box -33 -37 33 37
use M2M3_C_CDNS_7410113837434  M2M3_C_CDNS_7410113837434_13
timestamp 1748330293
transform 1 0 19366 0 1 34291
box -33 -37 33 37
use M2M3_C_CDNS_7410113837459  M2M3_C_CDNS_7410113837459_0
timestamp 1748330293
transform 1 0 20070 0 1 16293
box -33 -64 33 64
use M2M3_C_CDNS_7410113837459  M2M3_C_CDNS_7410113837459_1
timestamp 1748330293
transform 1 0 18058 0 1 34669
box -33 -64 33 64
use M2M3_C_CDNS_7410113837461  M2M3_C_CDNS_7410113837461_0
timestamp 1748330293
transform 1 0 17083 0 1 16913
box -50 -37 16 37
use M2M3_C_CDNS_7410113837461  M2M3_C_CDNS_7410113837461_1
timestamp 1748330293
transform 1 0 15071 0 1 35289
box -50 -37 16 37
use nfet_01v8_CDNS_741011383747  nfet_01v8_CDNS_741011383747_0
timestamp 1748330293
transform 1 0 14063 0 1 13972
box -71 -30 550 592
use nfet_01v8_CDNS_7410113837412  nfet_01v8_CDNS_7410113837412_0
timestamp 1748330293
transform 0 -1 9254 1 0 13547
box -239 -30 1079 192
use nfet_01v8_CDNS_7410113837412  nfet_01v8_CDNS_7410113837412_1
timestamp 1748330293
transform 0 -1 7242 1 0 31923
box -239 -30 1079 192
use nfet_01v8_CDNS_7410113837417  nfet_01v8_CDNS_7410113837417_0
timestamp 1748330293
transform 1 0 9885 0 1 12546
box -71 -154 109 2030
use nfet_01v8_CDNS_7410113837417  nfet_01v8_CDNS_7410113837417_1
timestamp 1748330293
transform 1 0 7873 0 1 30922
box -71 -154 109 2030
use nfet_01v8_CDNS_7410113837418  nfet_01v8_CDNS_7410113837418_0
timestamp 1748330293
transform -1 0 9657 0 1 12546
box -50 -154 101 2030
use nfet_01v8_CDNS_7410113837418  nfet_01v8_CDNS_7410113837418_1
timestamp 1748330293
transform -1 0 9829 0 1 12546
box -50 -154 101 2030
use nfet_01v8_CDNS_7410113837418  nfet_01v8_CDNS_7410113837418_2
timestamp 1748330293
transform -1 0 7645 0 1 30922
box -50 -154 101 2030
use nfet_01v8_CDNS_7410113837418  nfet_01v8_CDNS_7410113837418_3
timestamp 1748330293
transform -1 0 7817 0 1 30922
box -50 -154 101 2030
use nfet_01v8_CDNS_7410113837424  nfet_01v8_CDNS_7410113837424_0
timestamp 1748330293
transform 1 0 9713 0 1 12546
box -71 -154 80 2030
use nfet_01v8_CDNS_7410113837424  nfet_01v8_CDNS_7410113837424_1
timestamp 1748330293
transform 1 0 7701 0 1 30922
box -71 -154 80 2030
use nfet_01v8_CDNS_7410113837425  nfet_01v8_CDNS_7410113837425_0
timestamp 1748330293
transform 1 0 9541 0 1 12546
box -79 -154 80 2030
use nfet_01v8_CDNS_7410113837425  nfet_01v8_CDNS_7410113837425_1
timestamp 1748330293
transform 1 0 7529 0 1 30922
box -79 -154 80 2030
use nfet_01v8_CDNS_7410113837427  nfet_01v8_CDNS_7410113837427_0
timestamp 1748330293
transform 1 0 10219 0 1 14515
box -79 -154 80 230
use nfet_01v8_CDNS_7410113837427  nfet_01v8_CDNS_7410113837427_1
timestamp 1748330293
transform 1 0 8207 0 1 32891
box -79 -154 80 230
use nfet_01v8_CDNS_7410113837428  nfet_01v8_CDNS_7410113837428_0
timestamp 1748330293
transform 1 0 10291 0 1 14515
box -50 -154 109 230
use nfet_01v8_CDNS_7410113837428  nfet_01v8_CDNS_7410113837428_1
timestamp 1748330293
transform 1 0 8279 0 1 32891
box -50 -154 109 230
use nfet_01v8_CDNS_7410113837429  nfet_01v8_CDNS_7410113837429_0
timestamp 1748330293
transform 1 0 10513 0 1 14515
box -79 -154 109 230
use nfet_01v8_CDNS_7410113837429  nfet_01v8_CDNS_7410113837429_1
timestamp 1748330293
transform 1 0 11000 0 1 14515
box -79 -154 109 230
use nfet_01v8_CDNS_7410113837429  nfet_01v8_CDNS_7410113837429_2
timestamp 1748330293
transform 1 0 8501 0 1 32891
box -79 -154 109 230
use nfet_01v8_CDNS_7410113837429  nfet_01v8_CDNS_7410113837429_3
timestamp 1748330293
transform 1 0 8988 0 1 32891
box -79 -154 109 230
use nfet_01v8_CDNS_7410113837433  nfet_01v8_CDNS_7410113837433_0
timestamp 1748330293
transform -1 0 10823 0 1 14515
box -79 -154 80 230
use nfet_01v8_CDNS_7410113837433  nfet_01v8_CDNS_7410113837433_1
timestamp 1748330293
transform -1 0 8811 0 1 32891
box -79 -154 80 230
use nfet_01v8_CDNS_7410113837434  nfet_01v8_CDNS_7410113837434_0
timestamp 1748330293
transform 1 0 10707 0 1 14515
box -79 -154 101 230
use nfet_01v8_CDNS_7410113837434  nfet_01v8_CDNS_7410113837434_1
timestamp 1748330293
transform 1 0 8695 0 1 32891
box -79 -154 101 230
use nfet_01v8_CDNS_7410113837436  nfet_01v8_CDNS_7410113837436_0
timestamp 1748330293
transform -1 0 15781 0 1 13972
box -71 -30 579 592
use nfet_01v8_CDNS_7410113837436  nfet_01v8_CDNS_7410113837436_1
timestamp 1748330293
transform -1 0 17659 0 1 13972
box -71 -30 579 592
use nfet_01v8_CDNS_7410113837436  nfet_01v8_CDNS_7410113837436_2
timestamp 1748330293
transform -1 0 15647 0 1 32348
box -71 -30 579 592
use nfet_01v8_CDNS_7410113837437  nfet_01v8_CDNS_7410113837437_0
timestamp 1748330293
transform 1 0 15837 0 1 13972
box -50 -30 579 592
use nfet_01v8_CDNS_7410113837437  nfet_01v8_CDNS_7410113837437_1
timestamp 1748330293
transform 1 0 17715 0 1 13972
box -50 -30 579 592
use nfet_01v8_CDNS_7410113837437  nfet_01v8_CDNS_7410113837437_2
timestamp 1748330293
transform 1 0 15703 0 1 32348
box -50 -30 579 592
use nfet_01v8_CDNS_7410113837438  nfet_01v8_CDNS_7410113837438_0
timestamp 1748330293
transform 1 0 16497 0 1 13972
box -79 -30 579 592
use nfet_01v8_CDNS_7410113837438  nfet_01v8_CDNS_7410113837438_1
timestamp 1748330293
transform 1 0 14485 0 1 32348
box -79 -30 579 592
use nfet_01v8_CDNS_7410113837439  nfet_01v8_CDNS_7410113837439_0
timestamp 1748330293
transform 1 0 13507 0 1 13972
box -79 -30 550 592
use nfet_01v8_CDNS_7410113837440  nfet_01v8_CDNS_7410113837440_0
timestamp 1748330293
transform -1 0 15781 0 1 13418
box -71 -154 579 530
use nfet_01v8_CDNS_7410113837441  nfet_01v8_CDNS_7410113837441_0
timestamp 1748330293
transform -1 0 15119 0 1 13418
box -79 -154 571 530
use nfet_01v8_CDNS_7410113837442  nfet_01v8_CDNS_7410113837442_0
timestamp 1748330293
transform 1 0 13507 0 1 13418
box -79 -154 550 530
use nfet_01v8_CDNS_7410113837442  nfet_01v8_CDNS_7410113837442_1
timestamp 1748330293
transform -1 0 18215 0 1 13418
box -79 -154 550 530
use nfet_01v8_CDNS_7410113837442  nfet_01v8_CDNS_7410113837442_2
timestamp 1748330293
transform -1 0 16203 0 1 31794
box -79 -154 550 530
use nfet_01v8_CDNS_7410113837444  nfet_01v8_CDNS_7410113837444_0
timestamp 1748330293
transform -1 0 15119 0 1 13972
box -79 -30 571 592
use nfet_01v8_CDNS_7410113837446  nfet_01v8_CDNS_7410113837446_0
timestamp 1748330293
transform 1 0 16497 0 -1 13918
box -79 -30 579 654
use nfet_01v8_CDNS_7410113837446  nfet_01v8_CDNS_7410113837446_1
timestamp 1748330293
transform 1 0 14485 0 -1 32294
box -79 -30 579 654
use nfet_01v8_CDNS_7410113837447  nfet_01v8_CDNS_7410113837447_0
timestamp 1748330293
transform -1 0 17659 0 1 13418
box -71 -154 579 530
use nfet_01v8_CDNS_7410113837447  nfet_01v8_CDNS_7410113837447_1
timestamp 1748330293
transform -1 0 15647 0 1 31794
box -71 -154 579 530
use nfet_01v8_CDNS_7410113837448  nfet_01v8_CDNS_7410113837448_0
timestamp 1748330293
transform 1 0 14063 0 1 13418
box -71 -154 550 530
use nfet_01v8_CDNS_7410113837449  nfet_01v8_CDNS_7410113837449_0
timestamp 1748330293
transform 1 0 15837 0 1 13418
box -50 -154 579 530
use nfet_01v8_lvt_CDNS_741011383749  nfet_01v8_lvt_CDNS_741011383749_0
timestamp 1748330293
transform 1 0 12398 0 1 11304
box -37 -154 337 1492
use nfet_01v8_lvt_CDNS_7410113837416  nfet_01v8_lvt_CDNS_7410113837416_0
timestamp 1748330293
transform -1 0 12342 0 1 11304
box -71 -154 337 1492
use nfet_01v8_lvt_CDNS_7410113837435  nfet_01v8_lvt_CDNS_7410113837435_0
timestamp 1748330293
transform 1 0 21363 0 -1 15817
box -191 -30 109 230
use nfet_01v8_lvt_CDNS_7410113837435  nfet_01v8_lvt_CDNS_7410113837435_1
timestamp 1748330293
transform 1 0 19351 0 -1 34193
box -191 -30 109 230
use nfet_01v8_lvt_CDNS_7410113837445  nfet_01v8_lvt_CDNS_7410113837445_0
timestamp 1748330293
transform 1 0 12398 0 1 13018
box -71 -92 337 1554
use nfet_01v8_lvt_CDNS_7410113837452  nfet_01v8_lvt_CDNS_7410113837452_0
timestamp 1748330293
transform -1 0 13054 0 1 11304
box -79 -154 371 1492
use nfet_01v8_lvt_CDNS_7410113837452  nfet_01v8_lvt_CDNS_7410113837452_1
timestamp 1748330293
transform 1 0 11686 0 1 11304
box -79 -154 371 1492
use nfet_01v8_lvt_CDNS_7410113837454  nfet_01v8_lvt_CDNS_7410113837454_0
timestamp 1748330293
transform -1 0 13054 0 1 13018
box -79 -92 371 1554
use nfet_01v8_lvt_CDNS_7410113837455  nfet_01v8_lvt_CDNS_7410113837455_0
timestamp 1748330293
transform 1 0 11686 0 1 13018
box -79 -92 337 1554
use nfet_01v8_lvt_CDNS_7410113837456  nfet_01v8_lvt_CDNS_7410113837456_0
timestamp 1748330293
transform -1 0 12342 0 1 13018
box -37 -92 371 1554
use nfet_01v8_lvt_CDNS_7410113837474  nfet_01v8_lvt_CDNS_7410113837474_0
timestamp 1748330293
transform 0 -1 13734 1 0 12782
box -79 -30 221 230
use nfet_01v8_lvt_CDNS_7410113837474  nfet_01v8_lvt_CDNS_7410113837474_1
timestamp 1748330293
transform 0 -1 11722 1 0 31158
box -79 -30 221 230
use pfet_01v8_CDNS_7410113837410  pfet_01v8_CDNS_7410113837410_0
timestamp 1748330293
transform 0 -1 9814 -1 0 16022
box -236 -36 1089 202
use pfet_01v8_CDNS_7410113837410  pfet_01v8_CDNS_7410113837410_1
timestamp 1748330293
transform 0 -1 7802 -1 0 34398
box -236 -36 1089 202
use pfet_01v8_CDNS_7410113837413  pfet_01v8_CDNS_7410113837413_0
timestamp 1748330293
transform 1 0 16588 0 1 15055
box -50 -92 689 837
use pfet_01v8_CDNS_7410113837413  pfet_01v8_CDNS_7410113837413_1
timestamp 1748330293
transform 1 0 14576 0 1 33431
box -50 -92 689 837
use pfet_01v8_CDNS_7410113837414  pfet_01v8_CDNS_7410113837414_0
timestamp 1748330293
transform -1 0 16532 0 1 15055
box -81 -92 689 837
use pfet_01v8_CDNS_7410113837419  pfet_01v8_CDNS_7410113837419_0
timestamp 1748330293
transform -1 0 14476 0 1 15038
box -50 -92 281 872
use pfet_01v8_CDNS_7410113837420  pfet_01v8_CDNS_7410113837420_0
timestamp 1748330293
transform 0 -1 9574 -1 0 16022
box -236 -92 1089 146
use pfet_01v8_CDNS_7410113837420  pfet_01v8_CDNS_7410113837420_1
timestamp 1748330293
transform 0 -1 7562 -1 0 34398
box -236 -92 1089 146
use pfet_01v8_CDNS_7410113837421  pfet_01v8_CDNS_7410113837421_0
timestamp 1748330293
transform 1 0 10219 0 1 14847
box -89 -36 111 362
use pfet_01v8_CDNS_7410113837421  pfet_01v8_CDNS_7410113837421_1
timestamp 1748330293
transform 1 0 8207 0 1 33223
box -89 -36 111 362
use pfet_01v8_CDNS_7410113837422  pfet_01v8_CDNS_7410113837422_0
timestamp 1748330293
transform 1 0 11000 0 1 14847
box -89 -36 119 362
use pfet_01v8_CDNS_7410113837422  pfet_01v8_CDNS_7410113837422_1
timestamp 1748330293
transform 1 0 8501 0 1 33223
box -89 -36 119 362
use pfet_01v8_CDNS_7410113837422  pfet_01v8_CDNS_7410113837422_2
timestamp 1748330293
transform 1 0 10513 0 1 14847
box -89 -36 119 362
use pfet_01v8_CDNS_7410113837422  pfet_01v8_CDNS_7410113837422_3
timestamp 1748330293
transform 1 0 8988 0 1 33223
box -89 -36 119 362
use pfet_01v8_CDNS_7410113837423  pfet_01v8_CDNS_7410113837423_0
timestamp 1748330293
transform -1 0 10335 0 1 14847
box -89 -36 80 362
use pfet_01v8_CDNS_7410113837423  pfet_01v8_CDNS_7410113837423_1
timestamp 1748330293
transform -1 0 8323 0 1 33223
box -89 -36 80 362
use pfet_01v8_CDNS_7410113837426  pfet_01v8_CDNS_7410113837426_0
timestamp 1748330293
transform 0 -1 7342 -1 0 33428
box -201 -36 119 292
use pfet_01v8_CDNS_7410113837426  pfet_01v8_CDNS_7410113837426_1
timestamp 1748330293
transform 0 -1 9354 -1 0 15052
box -201 -36 119 292
use pfet_01v8_CDNS_7410113837430  pfet_01v8_CDNS_7410113837430_0
timestamp 1748330293
transform 1 0 17366 0 1 15055
box -89 -92 689 837
use pfet_01v8_CDNS_7410113837430  pfet_01v8_CDNS_7410113837430_1
timestamp 1748330293
transform -1 0 15754 0 1 15055
box -89 -92 689 837
use pfet_01v8_CDNS_7410113837430  pfet_01v8_CDNS_7410113837430_2
timestamp 1748330293
transform 1 0 15354 0 1 33431
box -89 -92 689 837
use pfet_01v8_CDNS_7410113837431  pfet_01v8_CDNS_7410113837431_0
timestamp 1748330293
transform 1 0 10793 0 1 14847
box -57 -36 119 362
use pfet_01v8_CDNS_7410113837431  pfet_01v8_CDNS_7410113837431_1
timestamp 1748330293
transform 1 0 8781 0 1 33223
box -57 -36 119 362
use pfet_01v8_CDNS_7410113837432  pfet_01v8_CDNS_7410113837432_0
timestamp 1748330293
transform 1 0 10721 0 1 14847
box -89 -36 87 362
use pfet_01v8_CDNS_7410113837432  pfet_01v8_CDNS_7410113837432_1
timestamp 1748330293
transform 1 0 8709 0 1 33223
box -89 -36 87 362
use pfet_01v8_CDNS_7410113837443  pfet_01v8_CDNS_7410113837443_0
timestamp 1748330293
transform -1 0 12906 0 1 15123
box -81 -92 289 636
use pfet_01v8_CDNS_7410113837443  pfet_01v8_CDNS_7410113837443_1
timestamp 1748330293
transform 1 0 12344 0 1 15123
box -81 -92 289 636
use pfet_01v8_CDNS_7410113837450  pfet_01v8_CDNS_7410113837450_0
timestamp 1748330293
transform 1 0 13708 0 1 16238
box -81 -92 650 1386
use pfet_01v8_CDNS_7410113837451  pfet_01v8_CDNS_7410113837451_0
timestamp 1748330293
transform -1 0 12032 0 1 15123
box -50 -92 401 692
use pfet_01v8_CDNS_7410113837451  pfet_01v8_CDNS_7410113837451_1
timestamp 1748330293
transform 1 0 13218 0 1 15123
box -50 -92 401 692
use pfet_01v8_CDNS_7410113837453  pfet_01v8_CDNS_7410113837453_0
timestamp 1748330293
transform -1 0 12288 0 1 15123
box -50 -92 281 692
use pfet_01v8_CDNS_7410113837453  pfet_01v8_CDNS_7410113837453_1
timestamp 1748330293
transform 1 0 12962 0 1 15123
box -50 -92 281 692
use pfet_01v8_CDNS_7410113837457  pfet_01v8_CDNS_7410113837457_0
timestamp 1748330293
transform 1 0 14532 0 1 15038
box -81 -92 289 872
use pfet_01v8_CDNS_7410113837458  pfet_01v8_CDNS_7410113837458_0
timestamp 1748330293
transform 1 0 14020 0 1 15038
box -89 -92 250 872
use pfet_01v8_CDNS_7410113837459  pfet_01v8_CDNS_7410113837459_0
timestamp 1748330293
transform 1 0 21800 0 1 16238
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837459  pfet_01v8_CDNS_7410113837459_1
timestamp 1748330293
transform 1 0 18786 0 1 16238
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837459  pfet_01v8_CDNS_7410113837459_2
timestamp 1748330293
transform 1 0 16774 0 1 34614
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837459  pfet_01v8_CDNS_7410113837459_3
timestamp 1748330293
transform 1 0 19788 0 1 34614
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837460  pfet_01v8_CDNS_7410113837460_0
timestamp 1748330293
transform 1 0 21800 0 1 17642
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837460  pfet_01v8_CDNS_7410113837460_1
timestamp 1748330293
transform 1 0 15020 0 1 17660
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837460  pfet_01v8_CDNS_7410113837460_2
timestamp 1748330293
transform -1 0 13652 0 1 17660
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837460  pfet_01v8_CDNS_7410113837460_3
timestamp 1748330293
transform -1 0 18730 0 1 17642
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837460  pfet_01v8_CDNS_7410113837460_4
timestamp 1748330293
transform -1 0 16718 0 1 36018
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_0
timestamp 1748330293
transform -1 0 21088 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_1
timestamp 1748330293
transform -1 0 12996 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_2
timestamp 1748330293
transform 1 0 15676 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_3
timestamp 1748330293
transform -1 0 18074 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_4
timestamp 1748330293
transform 1 0 19442 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_5
timestamp 1748330293
transform -1 0 16062 0 1 34614
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_6
timestamp 1748330293
transform 1 0 17430 0 1 34614
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837461  pfet_01v8_CDNS_7410113837461_7
timestamp 1748330293
transform -1 0 19076 0 1 34614
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_0
timestamp 1748330293
transform -1 0 21744 0 1 16238
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_1
timestamp 1748330293
transform 1 0 15020 0 1 16238
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_2
timestamp 1748330293
transform -1 0 13652 0 1 16238
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_3
timestamp 1748330293
transform -1 0 18730 0 1 16238
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_4
timestamp 1748330293
transform -1 0 16718 0 1 34614
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837462  pfet_01v8_CDNS_7410113837462_5
timestamp 1748330293
transform -1 0 19732 0 1 34614
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837463  pfet_01v8_CDNS_7410113837463_0
timestamp 1748330293
transform -1 0 24368 0 1 16238
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837463  pfet_01v8_CDNS_7410113837463_1
timestamp 1748330293
transform -1 0 22356 0 1 34614
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837464  pfet_01v8_CDNS_7410113837464_0
timestamp 1748330293
transform -1 0 17038 0 1 17660
box -89 -36 689 1512
use pfet_01v8_CDNS_7410113837464  pfet_01v8_CDNS_7410113837464_1
timestamp 1748330293
transform -1 0 12234 0 1 17660
box -89 -36 689 1512
use pfet_01v8_CDNS_7410113837464  pfet_01v8_CDNS_7410113837464_2
timestamp 1748330293
transform -1 0 15026 0 1 36036
box -89 -36 689 1512
use pfet_01v8_CDNS_7410113837465  pfet_01v8_CDNS_7410113837465_0
timestamp 1748330293
transform -1 0 14964 0 1 16238
box -81 -92 681 1386
use pfet_01v8_CDNS_7410113837466  pfet_01v8_CDNS_7410113837466_0
timestamp 1748330293
transform -1 0 14964 0 1 17660
box -81 -36 681 1512
use pfet_01v8_CDNS_7410113837467  pfet_01v8_CDNS_7410113837467_0
timestamp 1748330293
transform 1 0 13708 0 1 17660
box -81 -36 650 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_0
timestamp 1748330293
transform 1 0 25080 0 1 17642
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_1
timestamp 1748330293
transform -1 0 21088 0 1 17642
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_2
timestamp 1748330293
transform -1 0 12996 0 1 17660
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_3
timestamp 1748330293
transform 1 0 15676 0 1 17660
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_4
timestamp 1748330293
transform -1 0 18074 0 1 17642
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_5
timestamp 1748330293
transform 1 0 19442 0 1 17642
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_6
timestamp 1748330293
transform -1 0 16062 0 1 36018
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_7
timestamp 1748330293
transform 1 0 17430 0 1 36018
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_8
timestamp 1748330293
transform -1 0 19076 0 1 36018
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837468  pfet_01v8_CDNS_7410113837468_9
timestamp 1748330293
transform 1 0 23068 0 1 36018
box -50 -36 689 1512
use pfet_01v8_CDNS_7410113837469  pfet_01v8_CDNS_7410113837469_0
timestamp 1748330293
transform -1 0 12234 0 1 16238
box -89 -92 689 1386
use pfet_01v8_CDNS_7410113837469  pfet_01v8_CDNS_7410113837469_1
timestamp 1748330293
transform -1 0 17038 0 1 16238
box -89 -92 689 1386
use pfet_01v8_CDNS_7410113837469  pfet_01v8_CDNS_7410113837469_2
timestamp 1748330293
transform -1 0 15026 0 1 34614
box -89 -92 689 1386
use pfet_01v8_CDNS_7410113837470  pfet_01v8_CDNS_7410113837470_0
timestamp 1748330293
transform 1 0 23768 0 1 17642
box -81 -36 681 1512
use pfet_01v8_CDNS_7410113837470  pfet_01v8_CDNS_7410113837470_1
timestamp 1748330293
transform -1 0 21744 0 1 17642
box -81 -36 681 1512
use pfet_01v8_CDNS_7410113837470  pfet_01v8_CDNS_7410113837470_2
timestamp 1748330293
transform 1 0 18786 0 1 17642
box -81 -36 681 1512
use pfet_01v8_CDNS_7410113837470  pfet_01v8_CDNS_7410113837470_3
timestamp 1748330293
transform 1 0 16774 0 1 36018
box -81 -36 681 1512
use pfet_01v8_CDNS_7410113837471  pfet_01v8_CDNS_7410113837471_0
timestamp 1748330293
transform 1 0 24424 0 1 17642
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837472  pfet_01v8_CDNS_7410113837472_0
timestamp 1748330293
transform 1 0 25080 0 1 16238
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837472  pfet_01v8_CDNS_7410113837472_1
timestamp 1748330293
transform 1 0 23068 0 1 34614
box -50 -92 689 1386
use pfet_01v8_CDNS_7410113837473  pfet_01v8_CDNS_7410113837473_0
timestamp 1748330293
transform -1 0 23712 0 1 16238
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837473  pfet_01v8_CDNS_7410113837473_1
timestamp 1748330293
transform -1 0 21700 0 1 34614
box -50 -92 681 1386
use pfet_01v8_CDNS_7410113837475  pfet_01v8_CDNS_7410113837475_0
timestamp 1748330293
transform -1 0 25024 0 1 16238
box -81 -92 650 1386
use pfet_01v8_CDNS_7410113837475  pfet_01v8_CDNS_7410113837475_1
timestamp 1748330293
transform -1 0 23012 0 1 34614
box -81 -92 650 1386
use pfet_01v8_CDNS_7410113837476  pfet_01v8_CDNS_7410113837476_0
timestamp 1748330293
transform 1 0 22456 0 1 17642
box -50 -36 650 1512
use pfet_01v8_CDNS_7410113837477  pfet_01v8_CDNS_7410113837477_0
timestamp 1748330293
transform -1 0 23712 0 1 17642
box -50 -36 681 1512
use pfet_01v8_CDNS_7410113837478  pfet_01v8_CDNS_7410113837478_0
timestamp 1748330293
transform 1 0 22456 0 1 16238
box -50 -92 650 1386
use pfet_01v8_CDNS_7410113837478  pfet_01v8_CDNS_7410113837478_1
timestamp 1748330293
transform 1 0 20444 0 1 34614
box -50 -92 650 1386
use polyConn_CDNS_741011383740  polyConn_CDNS_741011383740_0
timestamp 1748330293
transform 1 0 21378 0 1 15915
box -26 -33 26 33
use polyConn_CDNS_741011383740  polyConn_CDNS_741011383740_1
timestamp 1748330293
transform 1 0 19366 0 1 34291
box -26 -33 26 33
use sky130_fd_pr__cap_mim_m3_1_WQ3WUD  sky130_fd_pr__cap_mim_m3_1_WQ3WUD_0
timestamp 1748330293
transform 1 0 18562 0 1 8608
box -2142 -3940 2142 3940
use sky130_fd_pr__cap_mim_m3_1_WQ3WUD  sky130_fd_pr__cap_mim_m3_1_WQ3WUD_1
timestamp 1748330293
transform 1 0 16550 0 1 26984
box -2142 -3940 2142 3940
use sky130_fd_pr__res_xhigh_po_0p35_VS6NPR  sky130_fd_pr__res_xhigh_po_0p35_VS6NPR_0
timestamp 1748330293
transform 0 1 15656 -1 0 12839
box -191 -1002 191 1002
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_0
timestamp 1748330293
transform 1 0 8659 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_1
timestamp 1748330293
transform 1 0 7763 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_2
timestamp 1748330293
transform 1 0 7651 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_3
timestamp 1748330293
transform 1 0 7875 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_4
timestamp 1748330293
transform 1 0 7987 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_5
timestamp 1748330293
transform 1 0 8099 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_6
timestamp 1748330293
transform 1 0 8211 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_7
timestamp 1748330293
transform 1 0 8323 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_8
timestamp 1748330293
transform 1 0 8435 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_9
timestamp 1748330293
transform 1 0 8547 0 1 15642
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_10
timestamp 1748330293
transform 1 0 6087 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_11
timestamp 1748330293
transform 1 0 6199 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_12
timestamp 1748330293
transform 1 0 6311 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_13
timestamp 1748330293
transform 1 0 5863 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_14
timestamp 1748330293
transform 1 0 5975 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_15
timestamp 1748330293
transform 1 0 5751 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_16
timestamp 1748330293
transform 1 0 5639 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_17
timestamp 1748330293
transform 1 0 6423 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_18
timestamp 1748330293
transform 1 0 6647 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_0p35_VXYPMA  sky130_fd_pr__res_xhigh_po_0p35_VXYPMA_19
timestamp 1748330293
transform 1 0 6535 0 1 34018
box -35 -2166 35 2166
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_0
timestamp 1748330293
transform 1 0 14729 0 1 8845
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_1
timestamp 1748330293
transform 1 0 14389 0 1 10285
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_2
timestamp 1748330293
transform 1 0 14729 0 1 10285
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_3
timestamp 1748330293
transform 1 0 14389 0 1 8845
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_4
timestamp 1748330293
transform 1 0 12377 0 1 27221
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_5
timestamp 1748330293
transform 1 0 12377 0 1 28661
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_6
timestamp 1748330293
transform 1 0 12717 0 1 27221
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_5RVTBE  sky130_fd_pr__res_xhigh_po_1p41_5RVTBE_7
timestamp 1748330293
transform 1 0 12717 0 1 28661
box -141 -645 141 645
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_0
timestamp 1748330293
transform 0 1 24824 -1 0 13161
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_1
timestamp 1748330293
transform 0 1 24824 -1 0 15141
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_2
timestamp 1748330293
transform 0 1 24824 -1 0 14811
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_3
timestamp 1748330293
transform 0 1 24824 -1 0 14481
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_4
timestamp 1748330293
transform 0 1 24824 -1 0 14149
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_5
timestamp 1748330293
transform 0 1 24824 -1 0 13821
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_6
timestamp 1748330293
transform 0 1 24824 -1 0 13491
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_B9H4MA  sky130_fd_pr__res_xhigh_po_1p41_B9H4MA_7
timestamp 1748330293
transform 0 1 24824 -1 0 12831
box -141 -976 141 976
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_0
timestamp 1748330293
transform 1 0 13639 0 1 10017
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_1
timestamp 1748330293
transform 1 0 15479 0 1 10017
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_2
timestamp 1748330293
transform 1 0 13639 0 1 4677
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_3
timestamp 1748330293
transform 1 0 13969 0 1 4677
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_4
timestamp 1748330293
transform 1 0 13969 0 1 10017
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_5
timestamp 1748330293
transform 1 0 15149 0 1 10017
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_6
timestamp 1748330293
transform 1 0 15479 0 1 4677
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_7
timestamp 1748330293
transform 1 0 15149 0 1 4677
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_8
timestamp 1748330293
transform 1 0 11627 0 1 28393
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_9
timestamp 1748330293
transform 1 0 11627 0 1 23053
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_10
timestamp 1748330293
transform 1 0 11957 0 1 28393
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_11
timestamp 1748330293
transform 1 0 11957 0 1 23053
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_12
timestamp 1748330293
transform 1 0 13137 0 1 28393
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_13
timestamp 1748330293
transform 1 0 13137 0 1 23053
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_14
timestamp 1748330293
transform 1 0 13467 0 1 28393
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_DHZREA  sky130_fd_pr__res_xhigh_po_1p41_DHZREA_15
timestamp 1748330293
transform 1 0 13467 0 1 23053
box -141 -2527 141 2527
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_0
timestamp 1748330293
transform 1 0 21371 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_1
timestamp 1748330293
transform 1 0 22019 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_2
timestamp 1748330293
transform 1 0 21695 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_3
timestamp 1748330293
transform 1 0 22343 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_4
timestamp 1748330293
transform 1 0 23639 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_5
timestamp 1748330293
transform 1 0 22667 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_6
timestamp 1748330293
transform 1 0 22991 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_7
timestamp 1748330293
transform 1 0 23315 0 1 14700
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_8
timestamp 1748330293
transform 1 0 20331 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_9
timestamp 1748330293
transform 1 0 20007 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_10
timestamp 1748330293
transform 1 0 19683 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_11
timestamp 1748330293
transform 1 0 19359 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_12
timestamp 1748330293
transform 1 0 21627 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_13
timestamp 1748330293
transform 1 0 21303 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_14
timestamp 1748330293
transform 1 0 20979 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_MV9HAT  sky130_fd_pr__res_xhigh_po_1p41_MV9HAT_15
timestamp 1748330293
transform 1 0 20655 0 1 33076
box -141 -652 141 652
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_0
timestamp 1748330293
transform -1 0 18645 0 -1 15163
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_1
timestamp 1748330293
transform -1 0 19295 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_2
timestamp 1748330293
transform -1 0 18647 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_3
timestamp 1748330293
transform -1 0 19293 0 -1 15163
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_4
timestamp 1748330293
transform -1 0 18971 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_5
timestamp 1748330293
transform -1 0 18969 0 -1 15163
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_6
timestamp 1748330293
transform -1 0 19943 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_7
timestamp 1748330293
transform -1 0 20267 0 -1 15137
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_8
timestamp 1748330293
transform -1 0 19619 0 -1 15137
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_9
timestamp 1748330293
transform -1 0 19943 0 -1 15137
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_10
timestamp 1748330293
transform -1 0 19619 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_11
timestamp 1748330293
transform -1 0 20591 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_12
timestamp 1748330293
transform -1 0 20591 0 -1 15137
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_13
timestamp 1748330293
transform -1 0 20915 0 -1 15137
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_14
timestamp 1748330293
transform -1 0 20267 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_15
timestamp 1748330293
transform -1 0 20915 0 -1 13715
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_16
timestamp 1748330293
transform -1 0 16631 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_17
timestamp 1748330293
transform -1 0 16631 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_18
timestamp 1748330293
transform -1 0 16955 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_19
timestamp 1748330293
transform -1 0 17279 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_20
timestamp 1748330293
transform -1 0 17279 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_21
timestamp 1748330293
transform -1 0 16955 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_22
timestamp 1748330293
transform -1 0 17603 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_23
timestamp 1748330293
transform -1 0 18575 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_24
timestamp 1748330293
transform -1 0 17603 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_25
timestamp 1748330293
transform -1 0 17927 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_26
timestamp 1748330293
transform -1 0 18575 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_27
timestamp 1748330293
transform -1 0 18251 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_28
timestamp 1748330293
transform -1 0 17927 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_29
timestamp 1748330293
transform -1 0 18251 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_30
timestamp 1748330293
transform -1 0 18899 0 -1 33607
box -141 -685 141 685
use sky130_fd_pr__res_xhigh_po_1p41_RG5DW9  sky130_fd_pr__res_xhigh_po_1p41_RG5DW9_31
timestamp 1748330293
transform -1 0 18899 0 -1 32195
box -141 -685 141 685
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0
array 0 2 1288 0 2 1288
timestamp 1748330293
transform 1 0 7156 0 1 24686
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
array 0 2 1288 0 2 1288
timestamp 1748330293
transform 1 0 9168 0 1 6310
box 0 0 1340 1340
<< labels >>
flabel metal4 s 27324 9690 27324 9690 0 FreeSans 7154 0 0 0 ua[0]
rlabel metal4 s 27324 9690 27324 9690 4 VDD
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 938 90 0 0 clk
port 2 nsew
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 938 90 0 0 ena
port 3 nsew
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 938 90 0 0 rst_n
port 4 nsew
flabel metal4 s 27234 0 27414 200 0 FreeSans 1876 0 0 0 ua[0]
port 5 nsew
flabel metal4 s 23370 0 23550 200 0 FreeSans 1876 0 0 0 ua[1]
port 6 nsew
flabel metal4 s 19506 0 19686 200 0 FreeSans 1876 0 0 0 ua[2]
port 7 nsew
flabel metal4 s 15642 0 15822 200 0 FreeSans 1876 0 0 0 ua[3]
port 8 nsew
flabel metal4 s 11778 0 11958 200 0 FreeSans 1876 0 0 0 ua[4]
port 9 nsew
flabel metal4 s 7914 0 8094 200 0 FreeSans 1876 0 0 0 ua[5]
port 10 nsew
flabel metal4 s 4050 0 4230 200 0 FreeSans 1876 0 0 0 ua[6]
port 11 nsew
flabel metal4 s 186 0 366 200 0 FreeSans 1876 0 0 0 ua[7]
port 12 nsew
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 938 90 0 0 ui_in[0]
port 13 nsew
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 938 90 0 0 ui_in[1]
port 14 nsew
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 938 90 0 0 ui_in[2]
port 15 nsew
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 938 90 0 0 ui_in[3]
port 16 nsew
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 938 90 0 0 ui_in[4]
port 17 nsew
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 938 90 0 0 ui_in[5]
port 18 nsew
rlabel metal4 s 23459 7330 23459 7330 4 VOUT
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 938 90 0 0 ui_in[6]
port 19 nsew
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 938 90 0 0 ui_in[7]
port 20 nsew
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 938 90 0 0 uio_in[0]
port 21 nsew
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 938 90 0 0 uio_in[1]
port 22 nsew
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 938 90 0 0 uio_in[2]
port 23 nsew
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 938 90 0 0 uio_in[3]
port 24 nsew
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 938 90 0 0 uio_in[4]
port 25 nsew
rlabel metal4 s 19596 1027 19596 1027 4 VDD_STRP
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 938 90 0 0 uio_in[5]
port 26 nsew
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 938 90 0 0 uio_in[6]
port 27 nsew
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 938 90 0 0 uio_in[7]
port 28 nsew
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 938 90 0 0 uio_oe[0]
port 29 nsew
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 938 90 0 0 uio_oe[1]
port 30 nsew
rlabel metal4 s 9546 17219 9546 17219 4 EN
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 938 90 0 0 uio_oe[2]
port 31 nsew
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 938 90 0 0 uio_oe[3]
port 32 nsew
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 938 90 0 0 uio_oe[4]
port 33 nsew
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 938 90 0 0 uio_oe[5]
port 34 nsew
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 938 90 0 0 uio_oe[6]
port 35 nsew
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 938 90 0 0 uio_oe[7]
port 36 nsew
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 938 90 0 0 uio_out[0]
port 37 nsew
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 938 90 0 0 uio_out[1]
port 38 nsew
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 938 90 0 0 uio_out[2]
port 39 nsew
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 938 90 0 0 uio_out[3]
port 40 nsew
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 938 90 0 0 uio_out[4]
port 41 nsew
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 938 90 0 0 uio_out[5]
port 42 nsew
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 938 90 0 0 uio_out[6]
port 43 nsew
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 938 90 0 0 uio_out[7]
port 44 nsew
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 938 90 0 0 uo_out[0]
port 45 nsew
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 938 90 0 0 uo_out[1]
port 46 nsew
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 938 90 0 0 uo_out[2]
port 47 nsew
rlabel metal4 s 7538 35538 7538 35538 4 EN1
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 938 90 0 0 uo_out[3]
port 48 nsew
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 938 90 0 0 uo_out[4]
port 49 nsew
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 938 90 0 0 uo_out[5]
port 50 nsew
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 938 90 0 0 uo_out[6]
port 51 nsew
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 938 90 0 0 uo_out[7]
port 52 nsew
flabel metal4 s 200 1000 440 44152 1 FreeSans 782 0 0 0 VDPWR
port 53 nsew
flabel metal4 s 800 1000 1040 44152 1 FreeSans 782 0 0 0 VGND
port 54 nsew
flabel metal4 s 1600 1000 1840 44152 1 FreeSans 782 0 0 0 VAPWR
port 55 nsew
rlabel metal2 s 25568 15234 25734 16900 4 VOUT
port 56 nsew
rlabel metal2 s 23556 33610 23722 35276 4 VOUT2
port 57 nsew
rlabel metal3 s 9022 34326 9088 34440 4 VDD2
port 58 nsew
rlabel metal3 s 8568 33666 8672 38340 4 EN_EXT1
port 59 nsew
rlabel metal1 s 8450 33493 8499 33547 4 VDD_STRP
port 60 nsew
rlabel metal1 s 10462 15117 10511 15171 4 VDD_STRP
port 60 nsew
rlabel metal1 s 9062 14752 9533 14804 4 EN
port 61 nsew
rlabel metal1 s 10618 15234 10652 15268 4 EN_EXT
port 62 nsew
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
