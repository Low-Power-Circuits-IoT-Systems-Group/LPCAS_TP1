magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 1304 -45 1350
rect -50 1270 -37 1304
rect -50 1236 -45 1270
rect -50 1202 -37 1236
rect -50 1168 -45 1202
rect -50 1134 -37 1168
rect -50 1100 -45 1134
rect -50 1066 -37 1100
rect -50 1032 -45 1066
rect -50 998 -37 1032
rect -50 964 -45 998
rect -50 930 -37 964
rect -50 896 -45 930
rect -50 862 -37 896
rect -50 828 -45 862
rect -50 794 -37 828
rect -50 760 -45 794
rect -50 726 -37 760
rect -50 692 -45 726
rect -50 658 -37 692
rect -50 624 -45 658
rect -50 590 -37 624
rect -50 556 -45 590
rect -50 522 -37 556
rect -50 488 -45 522
rect -50 454 -37 488
rect -50 420 -45 454
rect -50 386 -37 420
rect -50 352 -45 386
rect -50 318 -37 352
rect -50 284 -45 318
rect -50 250 -37 284
rect -50 216 -45 250
rect -50 182 -37 216
rect -50 148 -45 182
rect -50 114 -37 148
rect -50 80 -45 114
rect -50 46 -37 80
rect -50 0 -45 46
rect 611 0 650 1350
<< nwell >>
rect -81 -36 647 1512
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -45 1304 0 1350
rect -11 1270 0 1304
rect -45 1236 0 1270
rect -11 1202 0 1236
rect -45 1168 0 1202
rect -11 1134 0 1168
rect -45 1100 0 1134
rect -11 1066 0 1100
rect -45 1032 0 1066
rect -11 998 0 1032
rect -45 964 0 998
rect -11 930 0 964
rect -45 896 0 930
rect -11 862 0 896
rect -45 828 0 862
rect -11 794 0 828
rect -45 760 0 794
rect -11 726 0 760
rect -45 692 0 726
rect -11 658 0 692
rect -45 624 0 658
rect -11 590 0 624
rect -45 556 0 590
rect -11 522 0 556
rect -45 488 0 522
rect -11 454 0 488
rect -45 420 0 454
rect -11 386 0 420
rect -45 352 0 386
rect -11 318 0 352
rect -45 284 0 318
rect -11 250 0 284
rect -45 216 0 250
rect -11 182 0 216
rect -45 148 0 182
rect -11 114 0 148
rect -45 80 0 114
rect -11 46 0 80
rect -45 0 0 46
rect 600 0 611 1350
<< pdiffc >>
rect -45 1270 -11 1304
rect -45 1202 -11 1236
rect -45 1134 -11 1168
rect -45 1066 -11 1100
rect -45 998 -11 1032
rect -45 930 -11 964
rect -45 862 -11 896
rect -45 794 -11 828
rect -45 726 -11 760
rect -45 658 -11 692
rect -45 590 -11 624
rect -45 522 -11 556
rect -45 454 -11 488
rect -45 386 -11 420
rect -45 318 -11 352
rect -45 250 -11 284
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
<< nsubdiff >>
rect -45 1464 611 1476
rect -45 1430 -6 1464
rect 28 1430 62 1464
rect 96 1430 130 1464
rect 164 1430 198 1464
rect 232 1430 266 1464
rect 300 1430 334 1464
rect 368 1430 402 1464
rect 436 1430 470 1464
rect 504 1430 538 1464
rect 572 1430 611 1464
rect -45 1418 611 1430
<< nsubdiffcont >>
rect -6 1430 28 1464
rect 62 1430 96 1464
rect 130 1430 164 1464
rect 198 1430 232 1464
rect 266 1430 300 1464
rect 334 1430 368 1464
rect 402 1430 436 1464
rect 470 1430 504 1464
rect 538 1430 572 1464
<< poly >>
rect 0 1350 600 1380
rect 0 -30 600 0
<< locali >>
rect -43 1464 609 1474
rect -43 1430 -22 1464
rect 28 1430 50 1464
rect 96 1430 122 1464
rect 164 1430 194 1464
rect 232 1430 266 1464
rect 300 1430 334 1464
rect 372 1430 402 1464
rect 444 1430 470 1464
rect 516 1430 538 1464
rect 588 1430 609 1464
rect -43 1420 609 1430
rect -45 1304 -11 1350
rect -45 1236 -11 1270
rect -45 1168 -11 1202
rect -45 1100 -11 1134
rect -45 1032 -11 1066
rect -45 964 -11 998
rect -45 896 -11 930
rect -45 828 -11 862
rect -45 760 -11 794
rect -45 692 -11 726
rect -45 624 -11 658
rect -45 556 -11 590
rect -45 488 -11 522
rect -45 420 -11 454
rect -45 352 -11 386
rect -45 284 -11 318
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 0 -11 46
<< viali >>
rect -22 1430 -6 1464
rect -6 1430 12 1464
rect 50 1430 62 1464
rect 62 1430 84 1464
rect 122 1430 130 1464
rect 130 1430 156 1464
rect 194 1430 198 1464
rect 198 1430 228 1464
rect 266 1430 300 1464
rect 338 1430 368 1464
rect 368 1430 372 1464
rect 410 1430 436 1464
rect 436 1430 444 1464
rect 482 1430 504 1464
rect 504 1430 516 1464
rect 554 1430 572 1464
rect 572 1430 588 1464
<< metal1 >>
rect -43 1464 609 1474
rect -43 1430 -22 1464
rect 12 1430 50 1464
rect 84 1430 122 1464
rect 156 1430 194 1464
rect 228 1430 266 1464
rect 300 1430 338 1464
rect 372 1430 410 1464
rect 444 1430 482 1464
rect 516 1430 554 1464
rect 588 1430 609 1464
rect -43 1420 609 1430
<< end >>
