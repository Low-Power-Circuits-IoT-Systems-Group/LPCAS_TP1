magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< xpolycontact >>
rect -35 1734 35 2166
rect -35 -2166 35 -1734
<< xpolyres >>
rect -35 -1734 35 1734
<< viali >>
rect -17 2112 17 2146
rect -17 2040 17 2074
rect -17 1968 17 2002
rect -17 1896 17 1930
rect -17 1824 17 1858
rect -17 1752 17 1786
rect -17 -1787 17 -1753
rect -17 -1859 17 -1825
rect -17 -1931 17 -1897
rect -17 -2003 17 -1969
rect -17 -2075 17 -2041
rect -17 -2147 17 -2113
<< metal1 >>
rect -25 2146 25 2160
rect -25 2112 -17 2146
rect 17 2112 25 2146
rect -25 2074 25 2112
rect -25 2040 -17 2074
rect 17 2040 25 2074
rect -25 2002 25 2040
rect -25 1968 -17 2002
rect 17 1968 25 2002
rect -25 1930 25 1968
rect -25 1896 -17 1930
rect 17 1896 25 1930
rect -25 1858 25 1896
rect -25 1824 -17 1858
rect 17 1824 25 1858
rect -25 1786 25 1824
rect -25 1752 -17 1786
rect 17 1752 25 1786
rect -25 1739 25 1752
rect -25 -1753 25 -1739
rect -25 -1787 -17 -1753
rect 17 -1787 25 -1753
rect -25 -1825 25 -1787
rect -25 -1859 -17 -1825
rect 17 -1859 25 -1825
rect -25 -1897 25 -1859
rect -25 -1931 -17 -1897
rect 17 -1931 25 -1897
rect -25 -1969 25 -1931
rect -25 -2003 -17 -1969
rect 17 -2003 25 -1969
rect -25 -2041 25 -2003
rect -25 -2075 -17 -2041
rect 17 -2075 25 -2041
rect -25 -2113 25 -2075
rect -25 -2147 -17 -2113
rect 17 -2147 25 -2113
rect -25 -2160 25 -2147
<< end >>
