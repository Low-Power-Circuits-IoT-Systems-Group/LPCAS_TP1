magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -45 1329 -37 1363
rect -45 1261 -37 1295
rect -45 1193 -37 1227
rect -45 1125 -37 1159
rect -45 1057 -37 1091
rect -45 989 -37 1023
rect -45 921 -37 955
rect -45 853 -37 887
rect -45 785 -37 819
rect -45 717 -37 751
rect -45 649 -37 683
rect -45 581 -37 615
rect -45 513 -37 547
rect -45 445 -37 479
rect -45 377 -37 411
rect -45 309 -37 343
rect -45 241 -37 275
rect -45 173 -37 207
rect -45 105 -37 139
rect -45 37 -37 71
rect 311 0 330 1400
<< pwell >>
rect -71 -154 337 1426
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -45 1363 0 1400
rect -11 1329 0 1363
rect -45 1295 0 1329
rect -11 1261 0 1295
rect -45 1227 0 1261
rect -11 1193 0 1227
rect -45 1159 0 1193
rect -11 1125 0 1159
rect -45 1091 0 1125
rect -11 1057 0 1091
rect -45 1023 0 1057
rect -11 989 0 1023
rect -45 955 0 989
rect -11 921 0 955
rect -45 887 0 921
rect -11 853 0 887
rect -45 819 0 853
rect -11 785 0 819
rect -45 751 0 785
rect -11 717 0 751
rect -45 683 0 717
rect -11 649 0 683
rect -45 615 0 649
rect -11 581 0 615
rect -45 547 0 581
rect -11 513 0 547
rect -45 479 0 513
rect -11 445 0 479
rect -45 411 0 445
rect -11 377 0 411
rect -45 343 0 377
rect -11 309 0 343
rect -45 275 0 309
rect -11 241 0 275
rect -45 207 0 241
rect -11 173 0 207
rect -45 139 0 173
rect -11 105 0 139
rect -45 71 0 105
rect -11 37 0 71
rect -45 0 0 37
rect 300 0 311 1400
<< ndiffc >>
rect -45 1329 -11 1363
rect -45 1261 -11 1295
rect -45 1193 -11 1227
rect -45 1125 -11 1159
rect -45 1057 -11 1091
rect -45 989 -11 1023
rect -45 921 -11 955
rect -45 853 -11 887
rect -45 785 -11 819
rect -45 717 -11 751
rect -45 649 -11 683
rect -45 581 -11 615
rect -45 513 -11 547
rect -45 445 -11 479
rect -45 377 -11 411
rect -45 309 -11 343
rect -45 241 -11 275
rect -45 173 -11 207
rect -45 105 -11 139
rect -45 37 -11 71
<< psubdiff >>
rect -45 -82 311 -70
rect -45 -116 14 -82
rect 48 -116 82 -82
rect 116 -116 150 -82
rect 184 -116 218 -82
rect 252 -116 311 -82
rect -45 -128 311 -116
<< psubdiffcont >>
rect 14 -116 48 -82
rect 82 -116 116 -82
rect 150 -116 184 -82
rect 218 -116 252 -82
<< poly >>
rect 0 1482 300 1492
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1400 300 1448
rect 0 -30 300 0
<< polycont >>
rect 16 1448 50 1482
rect 94 1448 128 1482
rect 172 1448 206 1482
rect 250 1448 284 1482
<< locali >>
rect 0 1482 300 1488
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1442 300 1448
rect -45 1363 -11 1400
rect -45 1295 -11 1329
rect -45 1227 -11 1261
rect -45 1159 -11 1193
rect -45 1091 -11 1125
rect -45 1023 -11 1057
rect -45 955 -11 989
rect -45 887 -11 921
rect -45 819 -11 853
rect -45 751 -11 785
rect -45 683 -11 717
rect -45 615 -11 649
rect -45 547 -11 581
rect -45 479 -11 513
rect -45 411 -11 445
rect -45 343 -11 377
rect -45 275 -11 309
rect -45 207 -11 241
rect -45 139 -11 173
rect -45 71 -11 105
rect -45 0 -11 37
rect -43 -82 309 -72
rect -43 -116 8 -82
rect 48 -116 80 -82
rect 116 -116 150 -82
rect 186 -116 218 -82
rect 258 -116 309 -82
rect -43 -126 309 -116
<< viali >>
rect 16 1448 50 1482
rect 94 1448 128 1482
rect 172 1448 206 1482
rect 250 1448 284 1482
rect 8 -116 14 -82
rect 14 -116 42 -82
rect 80 -116 82 -82
rect 82 -116 114 -82
rect 152 -116 184 -82
rect 184 -116 186 -82
rect 224 -116 252 -82
rect 252 -116 258 -82
<< metal1 >>
rect 0 1482 300 1492
rect 0 1448 16 1482
rect 50 1448 94 1482
rect 128 1448 172 1482
rect 206 1448 250 1482
rect 284 1448 300 1482
rect 0 1438 300 1448
rect -43 -82 309 -72
rect -43 -116 8 -82
rect 42 -116 80 -82
rect 114 -116 152 -82
rect 186 -116 224 -82
rect 258 -116 309 -82
rect -43 -126 309 -116
<< end >>
