magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 675
<< nwell >>
rect -47 -36 689 837
<< pmos >>
rect 0 0 600 675
<< pdiff >>
rect -11 0 0 675
rect 600 626 653 675
rect 600 592 611 626
rect 645 592 653 626
rect 600 558 653 592
rect 600 524 611 558
rect 645 524 653 558
rect 600 490 653 524
rect 600 456 611 490
rect 645 456 653 490
rect 600 422 653 456
rect 600 388 611 422
rect 645 388 653 422
rect 600 354 653 388
rect 600 320 611 354
rect 645 320 653 354
rect 600 286 653 320
rect 600 252 611 286
rect 645 252 653 286
rect 600 218 653 252
rect 600 184 611 218
rect 645 184 653 218
rect 600 150 653 184
rect 600 116 611 150
rect 645 116 653 150
rect 600 82 653 116
rect 600 48 611 82
rect 645 48 653 82
rect 600 0 653 48
<< pdiffc >>
rect 611 592 645 626
rect 611 524 645 558
rect 611 456 645 490
rect 611 388 645 422
rect 611 320 645 354
rect 611 252 645 286
rect 611 184 645 218
rect 611 116 645 150
rect 611 48 645 82
<< nsubdiff >>
rect -11 789 653 801
rect -11 755 32 789
rect 66 755 100 789
rect 134 755 168 789
rect 202 755 236 789
rect 270 755 304 789
rect 338 755 372 789
rect 406 755 440 789
rect 474 755 508 789
rect 542 755 576 789
rect 610 755 653 789
rect -11 743 653 755
<< nsubdiffcont >>
rect 32 755 66 789
rect 100 755 134 789
rect 168 755 202 789
rect 236 755 270 789
rect 304 755 338 789
rect 372 755 406 789
rect 440 755 474 789
rect 508 755 542 789
rect 576 755 610 789
<< poly >>
rect 0 675 600 705
rect 0 -48 600 0
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< polycont >>
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< locali >>
rect -9 789 651 799
rect -9 755 16 789
rect 66 755 88 789
rect 134 755 160 789
rect 202 755 232 789
rect 270 755 304 789
rect 338 755 372 789
rect 410 755 440 789
rect 482 755 508 789
rect 554 755 576 789
rect 626 755 651 789
rect -9 745 651 755
rect 611 626 645 675
rect 611 558 645 592
rect 611 490 645 524
rect 611 422 645 456
rect 611 354 645 388
rect 611 286 645 320
rect 611 218 645 252
rect 611 150 645 184
rect 611 82 645 116
rect 611 0 645 48
rect 0 -48 600 -42
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -88 600 -82
<< viali >>
rect 16 755 32 789
rect 32 755 50 789
rect 88 755 100 789
rect 100 755 122 789
rect 160 755 168 789
rect 168 755 194 789
rect 232 755 236 789
rect 236 755 266 789
rect 304 755 338 789
rect 376 755 406 789
rect 406 755 410 789
rect 448 755 474 789
rect 474 755 482 789
rect 520 755 542 789
rect 542 755 554 789
rect 592 755 610 789
rect 610 755 626 789
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< metal1 >>
rect -9 789 651 799
rect -9 755 16 789
rect 50 755 88 789
rect 122 755 160 789
rect 194 755 232 789
rect 266 755 304 789
rect 338 755 376 789
rect 410 755 448 789
rect 482 755 520 789
rect 554 755 592 789
rect 626 755 651 789
rect -9 745 651 755
rect 0 -48 600 -38
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< end >>
