magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< nwell >>
rect -236 -36 1089 146
<< pmos >>
rect 0 0 1000 110
<< pdiff >>
rect -53 72 0 110
rect -53 38 -45 72
rect -11 38 0 72
rect -53 0 0 38
rect 1000 72 1053 110
rect 1000 38 1011 72
rect 1045 38 1053 72
rect 1000 0 1053 38
<< pdiffc >>
rect -45 38 -11 72
rect 1011 38 1045 72
<< nsubdiff >>
rect -200 72 -107 110
rect -200 38 -171 72
rect -137 38 -107 72
rect -200 0 -107 38
<< nsubdiffcont >>
rect -171 38 -137 72
<< poly >>
rect 0 192 1000 202
rect 0 158 16 192
rect 50 158 88 192
rect 122 158 160 192
rect 194 158 232 192
rect 266 158 304 192
rect 338 158 376 192
rect 410 158 448 192
rect 482 158 520 192
rect 554 158 592 192
rect 626 158 664 192
rect 698 158 736 192
rect 770 158 808 192
rect 842 158 879 192
rect 913 158 950 192
rect 984 158 1000 192
rect 0 110 1000 158
rect 0 -30 1000 0
<< polycont >>
rect 16 158 50 192
rect 88 158 122 192
rect 160 158 194 192
rect 232 158 266 192
rect 304 158 338 192
rect 376 158 410 192
rect 448 158 482 192
rect 520 158 554 192
rect 592 158 626 192
rect 664 158 698 192
rect 736 158 770 192
rect 808 158 842 192
rect 879 158 913 192
rect 950 158 984 192
<< locali >>
rect 0 192 1000 198
rect 0 158 16 192
rect 50 158 88 192
rect 128 158 160 192
rect 206 158 232 192
rect 284 158 304 192
rect 362 158 376 192
rect 440 158 448 192
rect 482 158 484 192
rect 518 158 520 192
rect 554 158 562 192
rect 626 158 640 192
rect 698 158 718 192
rect 770 158 796 192
rect 842 158 873 192
rect 913 158 950 192
rect 984 158 1000 192
rect 0 152 1000 158
rect -198 72 -109 110
rect -198 38 -171 72
rect -137 38 -109 72
rect -198 0 -109 38
rect -45 72 -11 110
rect -45 0 -11 38
rect 1011 72 1045 110
rect 1011 0 1045 38
<< viali >>
rect 16 158 50 192
rect 94 158 122 192
rect 122 158 128 192
rect 172 158 194 192
rect 194 158 206 192
rect 250 158 266 192
rect 266 158 284 192
rect 328 158 338 192
rect 338 158 362 192
rect 406 158 410 192
rect 410 158 440 192
rect 484 158 518 192
rect 562 158 592 192
rect 592 158 596 192
rect 640 158 664 192
rect 664 158 674 192
rect 718 158 736 192
rect 736 158 752 192
rect 796 158 808 192
rect 808 158 830 192
rect 873 158 879 192
rect 879 158 907 192
rect 950 158 984 192
rect -171 38 -137 72
<< metal1 >>
rect 0 192 1000 202
rect 0 158 16 192
rect 50 158 94 192
rect 128 158 172 192
rect 206 158 250 192
rect 284 158 328 192
rect 362 158 406 192
rect 440 158 484 192
rect 518 158 562 192
rect 596 158 640 192
rect 674 158 718 192
rect 752 158 796 192
rect 830 158 873 192
rect 907 158 950 192
rect 984 158 1000 192
rect 0 148 1000 158
rect -198 72 -109 110
rect -198 38 -171 72
rect -137 38 -109 72
rect -198 0 -109 38
<< end >>
