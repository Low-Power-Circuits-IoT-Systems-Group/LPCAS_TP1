magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 555 -45 600
rect -50 521 -37 555
rect -50 487 -45 521
rect -50 453 -37 487
rect -50 419 -45 453
rect -50 385 -37 419
rect -50 351 -45 385
rect -50 317 -37 351
rect -50 283 -45 317
rect -50 249 -37 283
rect -50 215 -45 249
rect -50 181 -37 215
rect -50 147 -45 181
rect -50 113 -37 147
rect -50 79 -45 113
rect -50 45 -37 79
rect -50 0 -45 45
<< nwell >>
rect -81 -36 289 636
<< pmos >>
rect 0 0 200 600
<< pdiff >>
rect -45 555 0 600
rect -11 521 0 555
rect -45 487 0 521
rect -11 453 0 487
rect -45 419 0 453
rect -11 385 0 419
rect -45 351 0 385
rect -11 317 0 351
rect -45 283 0 317
rect -11 249 0 283
rect -45 215 0 249
rect -11 181 0 215
rect -45 147 0 181
rect -11 113 0 147
rect -45 79 0 113
rect -11 45 0 79
rect -45 0 0 45
rect 200 555 253 600
rect 200 521 211 555
rect 245 521 253 555
rect 200 487 253 521
rect 200 453 211 487
rect 245 453 253 487
rect 200 419 253 453
rect 200 385 211 419
rect 245 385 253 419
rect 200 351 253 385
rect 200 317 211 351
rect 245 317 253 351
rect 200 283 253 317
rect 200 249 211 283
rect 245 249 253 283
rect 200 215 253 249
rect 200 181 211 215
rect 245 181 253 215
rect 200 147 253 181
rect 200 113 211 147
rect 245 113 253 147
rect 200 79 253 113
rect 200 45 211 79
rect 245 45 253 79
rect 200 0 253 45
<< pdiffc >>
rect -45 521 -11 555
rect -45 453 -11 487
rect -45 385 -11 419
rect -45 317 -11 351
rect -45 249 -11 283
rect -45 181 -11 215
rect -45 113 -11 147
rect -45 45 -11 79
rect 211 521 245 555
rect 211 453 245 487
rect 211 385 245 419
rect 211 317 245 351
rect 211 249 245 283
rect 211 181 245 215
rect 211 113 245 147
rect 211 45 245 79
<< poly >>
rect 0 600 200 630
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect -45 555 -11 600
rect -45 487 -11 521
rect -45 419 -11 453
rect -45 351 -11 385
rect -45 283 -11 317
rect -45 215 -11 249
rect -45 147 -11 181
rect -45 79 -11 113
rect -45 0 -11 45
rect 211 555 245 600
rect 211 487 245 521
rect 211 419 245 453
rect 211 351 245 385
rect 211 283 245 317
rect 211 215 245 249
rect 211 147 245 181
rect 211 79 245 113
rect 211 0 245 45
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
