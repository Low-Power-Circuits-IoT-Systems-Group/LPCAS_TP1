magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -34 -17 0 17
<< viali >>
rect -34 -17 0 17
<< metal1 >>
rect -43 17 9 32
rect -43 -17 -34 17
rect 0 -17 9 17
rect -43 -32 9 -17
<< end >>
