magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 77 200 79 362
rect 41 0 80 200
rect 77 -36 79 0
<< nwell >>
rect -89 -36 77 362
<< pmos >>
rect 0 0 30 200
<< pdiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 0 41 200
<< pdiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
<< nsubdiff >>
rect -53 314 41 326
rect -53 280 -23 314
rect 11 280 41 314
rect -53 268 41 280
<< nsubdiffcont >>
rect -23 280 11 314
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -51 314 39 324
rect -51 280 -23 314
rect 11 280 39 314
rect -51 270 39 280
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
<< viali >>
rect -23 280 11 314
<< metal1 >>
rect -51 314 39 324
rect -51 280 -23 314
rect 11 280 39 314
rect -51 270 39 280
<< end >>
