magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 545 471 550 500
rect 537 437 550 471
rect 545 403 550 437
rect 537 369 550 403
rect 545 335 550 369
rect 537 301 550 335
rect 545 267 550 301
rect 537 233 550 267
rect 545 199 550 233
rect 537 165 550 199
rect 545 131 550 165
rect 537 97 550 131
rect 545 63 550 97
rect 537 29 550 63
rect 545 0 550 29
<< pwell >>
rect -79 -154 571 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -53 471 0 500
rect -53 437 -45 471
rect -11 437 0 471
rect -53 403 0 437
rect -53 369 -45 403
rect -11 369 0 403
rect -53 335 0 369
rect -53 301 -45 335
rect -11 301 0 335
rect -53 267 0 301
rect -53 233 -45 267
rect -11 233 0 267
rect -53 199 0 233
rect -53 165 -45 199
rect -11 165 0 199
rect -53 131 0 165
rect -53 97 -45 131
rect -11 97 0 131
rect -53 63 0 97
rect -53 29 -45 63
rect -11 29 0 63
rect -53 0 0 29
rect 500 471 545 500
rect 500 437 511 471
rect 500 403 545 437
rect 500 369 511 403
rect 500 335 545 369
rect 500 301 511 335
rect 500 267 545 301
rect 500 233 511 267
rect 500 199 545 233
rect 500 165 511 199
rect 500 131 545 165
rect 500 97 511 131
rect 500 63 545 97
rect 500 29 511 63
rect 500 0 545 29
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< psubdiff >>
rect -53 -82 545 -70
rect -53 -116 -9 -82
rect 25 -116 59 -82
rect 93 -116 127 -82
rect 161 -116 195 -82
rect 229 -116 263 -82
rect 297 -116 331 -82
rect 365 -116 399 -82
rect 433 -116 467 -82
rect 501 -116 545 -82
rect -53 -128 545 -116
<< psubdiffcont >>
rect -9 -116 25 -82
rect 59 -116 93 -82
rect 127 -116 161 -82
rect 195 -116 229 -82
rect 263 -116 297 -82
rect 331 -116 365 -82
rect 399 -116 433 -82
rect 467 -116 501 -82
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
rect -51 -82 543 -72
rect -51 -116 -23 -82
rect 25 -116 49 -82
rect 93 -116 121 -82
rect 161 -116 193 -82
rect 229 -116 263 -82
rect 299 -116 331 -82
rect 371 -116 399 -82
rect 443 -116 467 -82
rect 515 -116 543 -82
rect -51 -126 543 -116
<< viali >>
rect -23 -116 -9 -82
rect -9 -116 11 -82
rect 49 -116 59 -82
rect 59 -116 83 -82
rect 121 -116 127 -82
rect 127 -116 155 -82
rect 193 -116 195 -82
rect 195 -116 227 -82
rect 265 -116 297 -82
rect 297 -116 299 -82
rect 337 -116 365 -82
rect 365 -116 371 -82
rect 409 -116 433 -82
rect 433 -116 443 -82
rect 481 -116 501 -82
rect 501 -116 515 -82
<< metal1 >>
rect -51 -82 543 -72
rect -51 -116 -23 -82
rect 11 -116 49 -82
rect 83 -116 121 -82
rect 155 -116 193 -82
rect 227 -116 265 -82
rect 299 -116 337 -82
rect 371 -116 409 -82
rect 443 -116 481 -82
rect 515 -116 543 -82
rect -51 -126 543 -116
<< end >>
