magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< pwell >>
rect -191 916 191 1002
rect -191 -916 -105 916
rect 105 -916 191 916
rect -191 -1002 191 -916
<< psubdiff >>
rect -165 942 -51 976
rect -17 942 17 976
rect 51 942 165 976
rect -165 867 -131 942
rect 131 867 165 942
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect -165 -942 -131 -867
rect 131 -942 165 -867
rect -165 -976 -51 -942
rect -17 -976 17 -942
rect 51 -976 165 -942
<< psubdiffcont >>
rect -51 942 -17 976
rect 17 942 51 976
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect -51 -976 -17 -942
rect 17 -976 51 -942
<< xpolycontact >>
rect -35 414 35 846
rect -35 -846 35 -414
<< xpolyres >>
rect -35 -414 35 414
<< locali >>
rect -165 942 -51 976
rect -17 942 17 976
rect 51 942 165 976
rect -165 867 -131 942
rect 131 867 165 942
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect -165 -942 -131 -867
rect 131 -942 165 -867
rect -165 -976 -51 -942
rect -17 -976 17 -942
rect 51 -976 165 -942
<< viali >>
rect -17 792 17 826
rect -17 720 17 754
rect -17 648 17 682
rect -17 576 17 610
rect -17 504 17 538
rect -17 432 17 466
rect -17 -467 17 -433
rect -17 -539 17 -505
rect -17 -611 17 -577
rect -17 -683 17 -649
rect -17 -755 17 -721
rect -17 -827 17 -793
<< metal1 >>
rect -25 826 25 840
rect -25 792 -17 826
rect 17 792 25 826
rect -25 754 25 792
rect -25 720 -17 754
rect 17 720 25 754
rect -25 682 25 720
rect -25 648 -17 682
rect 17 648 25 682
rect -25 610 25 648
rect -25 576 -17 610
rect 17 576 25 610
rect -25 538 25 576
rect -25 504 -17 538
rect 17 504 25 538
rect -25 466 25 504
rect -25 432 -17 466
rect 17 432 25 466
rect -25 419 25 432
rect -25 -433 25 -419
rect -25 -467 -17 -433
rect 17 -467 25 -433
rect -25 -505 25 -467
rect -25 -539 -17 -505
rect 17 -539 25 -505
rect -25 -577 25 -539
rect -25 -611 -17 -577
rect 17 -611 25 -577
rect -25 -649 25 -611
rect -25 -683 -17 -649
rect 17 -683 25 -649
rect -25 -721 25 -683
rect -25 -755 -17 -721
rect 17 -755 25 -721
rect -25 -793 25 -755
rect -25 -827 -17 -793
rect 17 -827 25 -793
rect -25 -840 25 -827
<< properties >>
string FIXED_BBOX -148 -959 148 959
<< end >>
