magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 500
<< pwell >>
rect -37 -26 579 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -11 0 0 500
rect 500 471 553 500
rect 500 437 511 471
rect 545 437 553 471
rect 500 403 553 437
rect 500 369 511 403
rect 545 369 553 403
rect 500 335 553 369
rect 500 301 511 335
rect 545 301 553 335
rect 500 267 553 301
rect 500 233 511 267
rect 545 233 553 267
rect 500 199 553 233
rect 500 165 511 199
rect 545 165 553 199
rect 500 131 553 165
rect 500 97 511 131
rect 545 97 553 131
rect 500 63 553 97
rect 500 29 511 63
rect 545 29 553 63
rect 500 0 553 29
<< ndiffc >>
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< poly >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 500 500 548
rect 0 -30 500 0
<< polycont >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< locali >>
rect 0 582 500 588
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 542 500 548
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
<< viali >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< metal1 >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 538 500 548
<< end >>
