magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 710
rect 245 678 250 710
rect 237 644 250 678
rect 245 610 250 644
rect 237 576 250 610
rect 245 542 250 576
rect 237 508 250 542
rect 245 474 250 508
rect 237 440 250 474
rect 245 406 250 440
rect 237 372 250 406
rect 245 338 250 372
rect 237 304 250 338
rect 245 270 250 304
rect 237 236 250 270
rect 245 202 250 236
rect 237 168 250 202
rect 245 134 250 168
rect 237 100 250 134
rect 245 66 250 100
rect 237 32 250 66
rect 245 0 250 32
<< nwell >>
rect -47 -36 281 872
<< pmos >>
rect 0 0 200 710
<< pdiff >>
rect -11 0 0 710
rect 200 678 245 710
rect 200 644 211 678
rect 200 610 245 644
rect 200 576 211 610
rect 200 542 245 576
rect 200 508 211 542
rect 200 474 245 508
rect 200 440 211 474
rect 200 406 245 440
rect 200 372 211 406
rect 200 338 245 372
rect 200 304 211 338
rect 200 270 245 304
rect 200 236 211 270
rect 200 202 245 236
rect 200 168 211 202
rect 200 134 245 168
rect 200 100 211 134
rect 200 66 245 100
rect 200 32 211 66
rect 200 0 245 32
<< pdiffc >>
rect 211 644 245 678
rect 211 576 245 610
rect 211 508 245 542
rect 211 440 245 474
rect 211 372 245 406
rect 211 304 245 338
rect 211 236 245 270
rect 211 168 245 202
rect 211 100 245 134
rect 211 32 245 66
<< nsubdiff >>
rect -11 824 245 836
rect -11 790 32 824
rect 66 790 100 824
rect 134 790 168 824
rect 202 790 245 824
rect -11 778 245 790
<< nsubdiffcont >>
rect 32 790 66 824
rect 100 790 134 824
rect 168 790 202 824
<< poly >>
rect 0 710 200 740
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect -9 824 243 834
rect -9 790 28 824
rect 66 790 100 824
rect 134 790 168 824
rect 206 790 243 824
rect -9 780 243 790
rect 211 678 245 710
rect 211 610 245 644
rect 211 542 245 576
rect 211 474 245 508
rect 211 406 245 440
rect 211 338 245 372
rect 211 270 245 304
rect 211 202 245 236
rect 211 134 245 168
rect 211 66 245 100
rect 211 0 245 32
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect 28 790 32 824
rect 32 790 62 824
rect 100 790 134 824
rect 172 790 202 824
rect 202 790 206 824
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect -9 824 243 834
rect -9 790 28 824
rect 62 790 100 824
rect 134 790 172 824
rect 206 790 243 824
rect -9 780 243 790
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
