magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -21 200
<< nwell >>
rect -57 -36 119 362
<< pmos >>
rect 0 0 30 200
<< pdiff >>
rect -21 0 0 200
rect 30 151 83 200
rect 30 117 41 151
rect 75 117 83 151
rect 30 83 83 117
rect 30 49 41 83
rect 75 49 83 83
rect 30 0 83 49
<< pdiffc >>
rect 41 117 75 151
rect 41 49 75 83
<< nsubdiff >>
rect -21 314 83 326
rect -21 280 14 314
rect 48 280 83 314
rect -21 268 83 280
<< nsubdiffcont >>
rect 14 280 48 314
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -19 314 81 324
rect -19 280 14 314
rect 48 280 81 314
rect -19 270 81 280
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
<< viali >>
rect 14 280 48 314
<< metal1 >>
rect -19 314 81 324
rect -19 280 14 314
rect 48 280 81 314
rect -19 270 81 280
<< end >>
