magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< pwell >>
rect -79 -26 221 226
<< nmoslvt >>
rect 0 0 30 200
<< ndiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 151 83 200
rect 30 117 41 151
rect 75 117 83 151
rect 30 83 83 117
rect 30 49 41 83
rect 75 49 83 83
rect 30 0 83 49
<< ndiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
rect 41 117 75 151
rect 41 49 75 83
<< psubdiff >>
rect 137 151 195 200
rect 137 117 149 151
rect 183 117 195 151
rect 137 83 195 117
rect 137 49 149 83
rect 183 49 195 83
rect 137 0 195 49
<< psubdiffcont >>
rect 149 117 183 151
rect 149 49 183 83
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
rect 139 153 193 200
rect 139 117 149 153
rect 183 117 193 153
rect 139 83 193 117
rect 139 47 149 83
rect 183 47 193 83
rect 139 0 193 47
<< viali >>
rect 149 151 183 153
rect 149 119 183 151
rect 149 49 183 81
rect 149 47 183 49
<< metal1 >>
rect 139 153 193 200
rect 139 119 149 153
rect 183 119 193 153
rect 139 81 193 119
rect 139 47 149 81
rect 183 47 193 81
rect 139 0 193 47
<< end >>
