magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 626 -45 675
rect -50 592 -37 626
rect -50 558 -45 592
rect -50 524 -37 558
rect -50 490 -45 524
rect -50 456 -37 490
rect -50 422 -45 456
rect -50 388 -37 422
rect -50 354 -45 388
rect -50 320 -37 354
rect -50 286 -45 320
rect -50 252 -37 286
rect -50 218 -45 252
rect -50 184 -37 218
rect -50 150 -45 184
rect -50 116 -37 150
rect -50 82 -45 116
rect -50 48 -37 82
rect -50 0 -45 48
<< nwell >>
rect -81 -36 689 837
<< pmos >>
rect 0 0 600 675
<< pdiff >>
rect -45 626 0 675
rect -11 592 0 626
rect -45 558 0 592
rect -11 524 0 558
rect -45 490 0 524
rect -11 456 0 490
rect -45 422 0 456
rect -11 388 0 422
rect -45 354 0 388
rect -11 320 0 354
rect -45 286 0 320
rect -11 252 0 286
rect -45 218 0 252
rect -11 184 0 218
rect -45 150 0 184
rect -11 116 0 150
rect -45 82 0 116
rect -11 48 0 82
rect -45 0 0 48
rect 600 626 653 675
rect 600 592 611 626
rect 645 592 653 626
rect 600 558 653 592
rect 600 524 611 558
rect 645 524 653 558
rect 600 490 653 524
rect 600 456 611 490
rect 645 456 653 490
rect 600 422 653 456
rect 600 388 611 422
rect 645 388 653 422
rect 600 354 653 388
rect 600 320 611 354
rect 645 320 653 354
rect 600 286 653 320
rect 600 252 611 286
rect 645 252 653 286
rect 600 218 653 252
rect 600 184 611 218
rect 645 184 653 218
rect 600 150 653 184
rect 600 116 611 150
rect 645 116 653 150
rect 600 82 653 116
rect 600 48 611 82
rect 645 48 653 82
rect 600 0 653 48
<< pdiffc >>
rect -45 592 -11 626
rect -45 524 -11 558
rect -45 456 -11 490
rect -45 388 -11 422
rect -45 320 -11 354
rect -45 252 -11 286
rect -45 184 -11 218
rect -45 116 -11 150
rect -45 48 -11 82
rect 611 592 645 626
rect 611 524 645 558
rect 611 456 645 490
rect 611 388 645 422
rect 611 320 645 354
rect 611 252 645 286
rect 611 184 645 218
rect 611 116 645 150
rect 611 48 645 82
<< nsubdiff >>
rect -45 789 653 801
rect -45 755 -19 789
rect 15 755 49 789
rect 83 755 117 789
rect 151 755 185 789
rect 219 755 253 789
rect 287 755 321 789
rect 355 755 389 789
rect 423 755 457 789
rect 491 755 525 789
rect 559 755 593 789
rect 627 755 653 789
rect -45 743 653 755
<< nsubdiffcont >>
rect -19 755 15 789
rect 49 755 83 789
rect 117 755 151 789
rect 185 755 219 789
rect 253 755 287 789
rect 321 755 355 789
rect 389 755 423 789
rect 457 755 491 789
rect 525 755 559 789
rect 593 755 627 789
<< poly >>
rect 0 675 600 705
rect 0 -48 600 0
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< polycont >>
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< locali >>
rect -43 789 651 799
rect -43 755 -19 789
rect 33 755 49 789
rect 105 755 117 789
rect 177 755 185 789
rect 249 755 253 789
rect 355 755 359 789
rect 423 755 431 789
rect 491 755 503 789
rect 559 755 575 789
rect 627 755 651 789
rect -43 745 651 755
rect -45 626 -11 675
rect -45 558 -11 592
rect -45 490 -11 524
rect -45 422 -11 456
rect -45 354 -11 388
rect -45 286 -11 320
rect -45 218 -11 252
rect -45 150 -11 184
rect -45 82 -11 116
rect -45 0 -11 48
rect 611 626 645 675
rect 611 558 645 592
rect 611 490 645 524
rect 611 422 645 456
rect 611 354 645 388
rect 611 286 645 320
rect 611 218 645 252
rect 611 150 645 184
rect 611 82 645 116
rect 611 0 645 48
rect 0 -48 600 -42
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -88 600 -82
<< viali >>
rect -1 755 15 789
rect 15 755 33 789
rect 71 755 83 789
rect 83 755 105 789
rect 143 755 151 789
rect 151 755 177 789
rect 215 755 219 789
rect 219 755 249 789
rect 287 755 321 789
rect 359 755 389 789
rect 389 755 393 789
rect 431 755 457 789
rect 457 755 465 789
rect 503 755 525 789
rect 525 755 537 789
rect 575 755 593 789
rect 593 755 609 789
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< metal1 >>
rect -43 789 651 799
rect -43 755 -1 789
rect 33 755 71 789
rect 105 755 143 789
rect 177 755 215 789
rect 249 755 287 789
rect 321 755 359 789
rect 393 755 431 789
rect 465 755 503 789
rect 537 755 575 789
rect 609 755 651 789
rect -43 745 651 755
rect 0 -48 600 -38
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< end >>
