magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 211 0 250 710
<< nwell >>
rect -89 -36 247 872
<< pmos >>
rect 0 0 200 710
<< pdiff >>
rect -53 678 0 710
rect -53 644 -45 678
rect -11 644 0 678
rect -53 610 0 644
rect -53 576 -45 610
rect -11 576 0 610
rect -53 542 0 576
rect -53 508 -45 542
rect -11 508 0 542
rect -53 474 0 508
rect -53 440 -45 474
rect -11 440 0 474
rect -53 406 0 440
rect -53 372 -45 406
rect -11 372 0 406
rect -53 338 0 372
rect -53 304 -45 338
rect -11 304 0 338
rect -53 270 0 304
rect -53 236 -45 270
rect -11 236 0 270
rect -53 202 0 236
rect -53 168 -45 202
rect -11 168 0 202
rect -53 134 0 168
rect -53 100 -45 134
rect -11 100 0 134
rect -53 66 0 100
rect -53 32 -45 66
rect -11 32 0 66
rect -53 0 0 32
rect 200 0 211 710
<< pdiffc >>
rect -45 644 -11 678
rect -45 576 -11 610
rect -45 508 -11 542
rect -45 440 -11 474
rect -45 372 -11 406
rect -45 304 -11 338
rect -45 236 -11 270
rect -45 168 -11 202
rect -45 100 -11 134
rect -45 32 -11 66
<< nsubdiff >>
rect -53 824 211 836
rect -53 790 -6 824
rect 28 790 62 824
rect 96 790 130 824
rect 164 790 211 824
rect -53 778 211 790
<< nsubdiffcont >>
rect -6 790 28 824
rect 62 790 96 824
rect 130 790 164 824
<< poly >>
rect 0 710 200 740
rect 0 -48 200 0
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< polycont >>
rect 16 -82 50 -48
rect 150 -82 184 -48
<< locali >>
rect -51 824 209 834
rect -51 790 -10 824
rect 28 790 62 824
rect 96 790 130 824
rect 168 790 209 824
rect -51 780 209 790
rect -45 678 -11 710
rect -45 610 -11 644
rect -45 542 -11 576
rect -45 474 -11 508
rect -45 406 -11 440
rect -45 338 -11 372
rect -45 270 -11 304
rect -45 202 -11 236
rect -45 134 -11 168
rect -45 66 -11 100
rect -45 0 -11 32
rect 0 -48 200 -42
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -88 200 -82
<< viali >>
rect -10 790 -6 824
rect -6 790 24 824
rect 62 790 96 824
rect 134 790 164 824
rect 164 790 168 824
rect 16 -82 50 -48
rect 150 -82 184 -48
<< metal1 >>
rect -51 824 209 834
rect -51 790 -10 824
rect 24 790 62 824
rect 96 790 134 824
rect 168 790 209 824
rect -51 780 209 790
rect 0 -48 200 -38
rect 0 -82 16 -48
rect 50 -82 150 -48
rect 184 -82 200 -48
rect 0 -92 200 -82
<< end >>
