magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< xpolycontact >>
rect -141 2095 141 2527
rect -141 -2527 141 -2095
<< xpolyres >>
rect -141 -2095 141 2095
<< viali >>
rect -125 2113 125 2507
rect -125 -2508 125 -2114
<< metal1 >>
rect -131 2507 131 2521
rect -131 2113 -125 2507
rect 125 2113 131 2507
rect -131 2100 131 2113
rect -131 -2114 131 -2100
rect -131 -2508 -125 -2114
rect 125 -2508 131 -2114
rect -131 -2521 131 -2508
<< end >>
