magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -26 90 26 101
rect -26 26 26 38
rect -26 -38 26 -26
rect -26 -101 26 -90
<< via1 >>
rect -26 38 26 90
rect -26 -26 26 26
rect -26 -90 26 -38
<< metal2 >>
rect -32 38 -26 90
rect 26 38 32 90
rect -32 26 32 38
rect -32 -26 -26 26
rect 26 -26 32 26
rect -32 -38 32 -26
rect -32 -90 -26 -38
rect 26 -90 32 -38
<< end >>
