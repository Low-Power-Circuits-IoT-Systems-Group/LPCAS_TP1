VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_LPCAS_TP1
  CLASS BLOCK ;
  FOREIGN tt_um_LPCAS_TP1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN VDD
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 96.900 ;
    END
    PORT
      LAYER li1 ;
        RECT 57.285 77.470 57.455 77.640 ;
    END
    PORT
      LAYER li1 ;
        RECT 47.225 169.350 47.395 169.520 ;
    END
  END VDD
  PIN ua[1]
    ANTENNAGATEAREA 18.150000 ;
    ANTENNADIFFAREA 15.650000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNADIFFAREA 7.542800 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 7.500000 ;
    ANTENNADIFFAREA 10.934999 ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN GND
    ANTENNAGATEAREA 481.120178 ;
    ANTENNADIFFAREA 457.449188 ;
    PORT
      LAYER li1 ;
        RECT 50.420 71.930 57.230 72.230 ;
    END
    PORT
      LAYER li1 ;
        RECT 40.360 163.810 47.170 164.110 ;
    END
  END GND
  PIN ui_in[1]
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN VOUT
    ANTENNAGATEAREA 18.150000 ;
    ANTENNADIFFAREA 15.650000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.740 73.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 127.840 76.170 128.670 84.500 ;
    END
  END VOUT
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN VDD2
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met3 ;
        RECT 45.110 171.630 45.440 172.200 ;
    END
  END VDD2
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN VDD_STRP
    ANTENNADIFFAREA 7.542800 ;
    PORT
      LAYER met4 ;
        RECT 97.540 0.000 98.420 10.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.310 75.585 52.555 75.855 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.250 167.465 42.495 167.735 ;
    END
  END VDD_STRP
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN EN
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 47.480 74.060 47.980 98.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 45.310 73.760 47.665 74.020 ;
    END
  END EN
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN EN_EXT
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met1 ;
        RECT 53.090 76.170 53.260 76.340 ;
    END
  END EN_EXT
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN VOUT2
    ANTENNAGATEAREA 7.500000 ;
    ANTENNADIFFAREA 10.934999 ;
    PORT
      LAYER met2 ;
        RECT 117.780 168.050 118.610 176.380 ;
    END
  END VOUT2
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN EN1
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 37.400 166.020 37.980 189.360 ;
    END
  END EN1
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN EN_EXT1
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met3 ;
        RECT 42.840 168.330 43.360 191.700 ;
    END
  END EN_EXT1
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.200 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    ANTENNADIFFAREA 7.542800 ;
    PORT
      LAYER met4 ;
        RECT 8.000 5.000 9.200 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 34.140 31.550 129.515 188.360 ;
      LAYER li1 ;
        RECT 28.020 169.690 129.335 188.180 ;
        RECT 28.020 169.180 47.055 169.690 ;
        RECT 47.565 169.180 129.335 169.690 ;
        RECT 28.020 164.280 129.335 169.180 ;
        RECT 28.020 163.640 40.190 164.280 ;
        RECT 47.340 163.640 129.335 164.280 ;
        RECT 28.020 77.810 129.335 163.640 ;
        RECT 28.020 77.300 57.115 77.810 ;
        RECT 57.625 77.300 129.335 77.810 ;
        RECT 28.020 72.400 129.335 77.300 ;
        RECT 28.020 71.760 50.250 72.400 ;
        RECT 57.400 71.760 129.335 72.400 ;
        RECT 28.020 10.750 129.335 71.760 ;
      LAYER met1 ;
        RECT 28.030 168.015 129.010 187.550 ;
        RECT 28.030 167.185 41.970 168.015 ;
        RECT 42.775 167.185 129.010 168.015 ;
        RECT 28.030 76.620 129.010 167.185 ;
        RECT 28.030 76.135 52.810 76.620 ;
        RECT 28.030 75.305 52.030 76.135 ;
        RECT 53.540 75.890 129.010 76.620 ;
        RECT 52.835 75.305 129.010 75.890 ;
        RECT 28.030 74.300 129.010 75.305 ;
        RECT 28.030 73.480 45.030 74.300 ;
        RECT 47.945 73.480 129.010 74.300 ;
        RECT 28.030 10.750 129.010 73.480 ;
      LAYER met2 ;
        RECT 27.980 176.660 129.060 180.100 ;
        RECT 27.980 167.770 117.500 176.660 ;
        RECT 118.890 167.770 129.060 176.660 ;
        RECT 27.980 84.780 129.060 167.770 ;
        RECT 27.980 75.890 127.560 84.780 ;
        RECT 128.950 75.890 129.060 84.780 ;
        RECT 27.980 33.890 129.060 75.890 ;
      LAYER met3 ;
        RECT 3.990 192.100 129.070 192.320 ;
        RECT 3.990 167.930 42.440 192.100 ;
        RECT 43.760 172.600 129.070 192.100 ;
        RECT 43.760 171.230 44.710 172.600 ;
        RECT 45.840 171.230 129.070 172.600 ;
        RECT 43.760 167.930 129.070 171.230 ;
        RECT 3.990 23.940 129.070 167.930 ;
      LAYER met4 ;
        RECT 9.200 224.360 14.630 224.760 ;
        RECT 15.730 224.360 17.390 224.760 ;
        RECT 18.490 224.360 20.150 224.760 ;
        RECT 21.250 224.360 22.910 224.760 ;
        RECT 24.010 224.360 25.670 224.760 ;
        RECT 26.770 224.360 28.430 224.760 ;
        RECT 29.530 224.360 31.190 224.760 ;
        RECT 32.290 224.360 33.950 224.760 ;
        RECT 35.050 224.360 36.710 224.760 ;
        RECT 37.810 224.360 39.470 224.760 ;
        RECT 40.570 224.360 42.230 224.760 ;
        RECT 43.330 224.360 44.990 224.760 ;
        RECT 46.090 224.360 47.750 224.760 ;
        RECT 48.850 224.360 50.510 224.760 ;
        RECT 51.610 224.360 53.270 224.760 ;
        RECT 54.370 224.360 56.030 224.760 ;
        RECT 57.130 224.360 58.790 224.760 ;
        RECT 59.890 224.360 61.550 224.760 ;
        RECT 62.650 224.360 64.310 224.760 ;
        RECT 65.410 224.360 67.070 224.760 ;
        RECT 68.170 224.360 69.830 224.760 ;
        RECT 70.930 224.360 72.590 224.760 ;
        RECT 73.690 224.360 75.350 224.760 ;
        RECT 76.450 224.360 78.110 224.760 ;
        RECT 79.210 224.360 80.870 224.760 ;
        RECT 81.970 224.360 83.630 224.760 ;
        RECT 84.730 224.360 86.390 224.760 ;
        RECT 87.490 224.360 89.150 224.760 ;
        RECT 90.250 224.360 91.910 224.760 ;
        RECT 93.010 224.360 94.670 224.760 ;
        RECT 95.770 224.360 97.430 224.760 ;
        RECT 98.530 224.360 100.190 224.760 ;
        RECT 101.290 224.360 102.950 224.760 ;
        RECT 104.050 224.360 105.710 224.760 ;
        RECT 106.810 224.360 108.470 224.760 ;
        RECT 109.570 224.360 111.230 224.760 ;
        RECT 112.330 224.360 113.990 224.760 ;
        RECT 115.090 224.360 116.750 224.760 ;
        RECT 117.850 224.360 119.510 224.760 ;
        RECT 120.610 224.360 122.270 224.760 ;
        RECT 123.370 224.360 125.030 224.760 ;
        RECT 126.130 224.360 127.790 224.760 ;
        RECT 128.890 224.360 130.550 224.760 ;
        RECT 131.650 224.360 136.170 224.760 ;
        RECT 9.200 221.160 136.170 224.360 ;
        RECT 9.600 189.760 136.170 221.160 ;
        RECT 9.600 165.620 37.000 189.760 ;
        RECT 38.380 165.620 136.170 189.760 ;
        RECT 9.600 98.530 136.170 165.620 ;
        RECT 9.600 73.660 47.080 98.530 ;
        RECT 48.380 97.300 136.170 98.530 ;
        RECT 48.380 73.700 135.770 97.300 ;
        RECT 48.380 73.660 116.450 73.700 ;
        RECT 9.600 10.670 116.450 73.660 ;
        RECT 9.600 4.600 97.140 10.670 ;
        RECT 9.200 1.400 97.140 4.600 ;
        RECT 98.820 1.400 116.450 10.670 ;
        RECT 118.140 1.400 135.770 73.700 ;
        RECT 9.200 1.000 19.850 1.400 ;
        RECT 21.550 1.000 39.170 1.400 ;
        RECT 40.870 1.000 58.490 1.400 ;
        RECT 60.190 1.000 77.810 1.400 ;
        RECT 79.510 1.000 97.130 1.400 ;
        RECT 98.830 1.000 116.450 1.400 ;
        RECT 118.150 1.000 135.770 1.400 ;
  END
END tt_um_LPCAS_TP1
END LIBRARY

