magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -26 314 26 353
rect -26 250 26 262
rect -26 186 26 198
rect -26 122 26 134
rect -26 58 26 70
rect -26 -6 26 6
rect -26 -70 26 -58
rect -26 -134 26 -122
rect -26 -198 26 -186
rect -26 -262 26 -250
rect -26 -353 26 -314
<< via1 >>
rect -26 262 26 314
rect -26 198 26 250
rect -26 134 26 186
rect -26 70 26 122
rect -26 6 26 58
rect -26 -58 26 -6
rect -26 -122 26 -70
rect -26 -186 26 -134
rect -26 -250 26 -198
rect -26 -314 26 -262
<< metal2 >>
rect -26 314 26 320
rect -26 250 26 262
rect -26 186 26 198
rect -26 122 26 134
rect -26 58 26 70
rect -26 -6 26 6
rect -26 -70 26 -58
rect -26 -134 26 -122
rect -26 -198 26 -186
rect -26 -262 26 -250
rect -26 -320 26 -314
<< end >>
