magic
tech sky130A
timestamp 1741700111
<< metal1 >>
rect -48 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 48 13
<< via1 >>
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
<< metal2 >>
rect -48 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 48 13
<< end >>
