magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -11 1350
<< nwell >>
rect -47 -36 689 1512
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -11 0 0 1350
rect 600 1304 653 1350
rect 600 1270 611 1304
rect 645 1270 653 1304
rect 600 1236 653 1270
rect 600 1202 611 1236
rect 645 1202 653 1236
rect 600 1168 653 1202
rect 600 1134 611 1168
rect 645 1134 653 1168
rect 600 1100 653 1134
rect 600 1066 611 1100
rect 645 1066 653 1100
rect 600 1032 653 1066
rect 600 998 611 1032
rect 645 998 653 1032
rect 600 964 653 998
rect 600 930 611 964
rect 645 930 653 964
rect 600 896 653 930
rect 600 862 611 896
rect 645 862 653 896
rect 600 828 653 862
rect 600 794 611 828
rect 645 794 653 828
rect 600 760 653 794
rect 600 726 611 760
rect 645 726 653 760
rect 600 692 653 726
rect 600 658 611 692
rect 645 658 653 692
rect 600 624 653 658
rect 600 590 611 624
rect 645 590 653 624
rect 600 556 653 590
rect 600 522 611 556
rect 645 522 653 556
rect 600 488 653 522
rect 600 454 611 488
rect 645 454 653 488
rect 600 420 653 454
rect 600 386 611 420
rect 645 386 653 420
rect 600 352 653 386
rect 600 318 611 352
rect 645 318 653 352
rect 600 284 653 318
rect 600 250 611 284
rect 645 250 653 284
rect 600 216 653 250
rect 600 182 611 216
rect 645 182 653 216
rect 600 148 653 182
rect 600 114 611 148
rect 645 114 653 148
rect 600 80 653 114
rect 600 46 611 80
rect 645 46 653 80
rect 600 0 653 46
<< pdiffc >>
rect 611 1270 645 1304
rect 611 1202 645 1236
rect 611 1134 645 1168
rect 611 1066 645 1100
rect 611 998 645 1032
rect 611 930 645 964
rect 611 862 645 896
rect 611 794 645 828
rect 611 726 645 760
rect 611 658 645 692
rect 611 590 645 624
rect 611 522 645 556
rect 611 454 645 488
rect 611 386 645 420
rect 611 318 645 352
rect 611 250 645 284
rect 611 182 645 216
rect 611 114 645 148
rect 611 46 645 80
<< nsubdiff >>
rect -11 1464 653 1476
rect -11 1430 32 1464
rect 66 1430 100 1464
rect 134 1430 168 1464
rect 202 1430 236 1464
rect 270 1430 304 1464
rect 338 1430 372 1464
rect 406 1430 440 1464
rect 474 1430 508 1464
rect 542 1430 576 1464
rect 610 1430 653 1464
rect -11 1418 653 1430
<< nsubdiffcont >>
rect 32 1430 66 1464
rect 100 1430 134 1464
rect 168 1430 202 1464
rect 236 1430 270 1464
rect 304 1430 338 1464
rect 372 1430 406 1464
rect 440 1430 474 1464
rect 508 1430 542 1464
rect 576 1430 610 1464
<< poly >>
rect 0 1350 600 1380
rect 0 -30 600 0
<< locali >>
rect -9 1464 651 1474
rect -9 1430 16 1464
rect 66 1430 88 1464
rect 134 1430 160 1464
rect 202 1430 232 1464
rect 270 1430 304 1464
rect 338 1430 372 1464
rect 410 1430 440 1464
rect 482 1430 508 1464
rect 554 1430 576 1464
rect 626 1430 651 1464
rect -9 1420 651 1430
rect 611 1304 645 1350
rect 611 1236 645 1270
rect 611 1168 645 1202
rect 611 1100 645 1134
rect 611 1032 645 1066
rect 611 964 645 998
rect 611 896 645 930
rect 611 828 645 862
rect 611 760 645 794
rect 611 692 645 726
rect 611 624 645 658
rect 611 556 645 590
rect 611 488 645 522
rect 611 420 645 454
rect 611 352 645 386
rect 611 284 645 318
rect 611 216 645 250
rect 611 148 645 182
rect 611 80 645 114
rect 611 0 645 46
<< viali >>
rect 16 1430 32 1464
rect 32 1430 50 1464
rect 88 1430 100 1464
rect 100 1430 122 1464
rect 160 1430 168 1464
rect 168 1430 194 1464
rect 232 1430 236 1464
rect 236 1430 266 1464
rect 304 1430 338 1464
rect 376 1430 406 1464
rect 406 1430 410 1464
rect 448 1430 474 1464
rect 474 1430 482 1464
rect 520 1430 542 1464
rect 542 1430 554 1464
rect 592 1430 610 1464
rect 610 1430 626 1464
<< metal1 >>
rect -9 1464 651 1474
rect -9 1430 16 1464
rect 50 1430 88 1464
rect 122 1430 160 1464
rect 194 1430 232 1464
rect 266 1430 304 1464
rect 338 1430 376 1464
rect 410 1430 448 1464
rect 482 1430 520 1464
rect 554 1430 592 1464
rect 626 1430 651 1464
rect -9 1420 651 1430
<< end >>
