magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 1304 -45 1350
rect 645 1304 650 1350
rect -50 1270 -37 1304
rect 637 1270 650 1304
rect -50 1236 -45 1270
rect 645 1236 650 1270
rect -50 1202 -37 1236
rect 637 1202 650 1236
rect -50 1168 -45 1202
rect 645 1168 650 1202
rect -50 1134 -37 1168
rect 637 1134 650 1168
rect -50 1100 -45 1134
rect 645 1100 650 1134
rect -50 1066 -37 1100
rect 637 1066 650 1100
rect -50 1032 -45 1066
rect 645 1032 650 1066
rect -50 998 -37 1032
rect 637 998 650 1032
rect -50 964 -45 998
rect 645 964 650 998
rect -50 930 -37 964
rect 637 930 650 964
rect -50 896 -45 930
rect 645 896 650 930
rect -50 862 -37 896
rect 637 862 650 896
rect -50 828 -45 862
rect 645 828 650 862
rect -50 794 -37 828
rect 637 794 650 828
rect -50 760 -45 794
rect 645 760 650 794
rect -50 726 -37 760
rect 637 726 650 760
rect -50 692 -45 726
rect 645 692 650 726
rect -50 658 -37 692
rect 637 658 650 692
rect -50 624 -45 658
rect 645 624 650 658
rect -50 590 -37 624
rect 637 590 650 624
rect -50 556 -45 590
rect 645 556 650 590
rect -50 522 -37 556
rect 637 522 650 556
rect -50 488 -45 522
rect 645 488 650 522
rect -50 454 -37 488
rect 637 454 650 488
rect -50 420 -45 454
rect 645 420 650 454
rect -50 386 -37 420
rect 637 386 650 420
rect -50 352 -45 386
rect 645 352 650 386
rect -50 318 -37 352
rect 637 318 650 352
rect -50 284 -45 318
rect 645 284 650 318
rect -50 250 -37 284
rect 637 250 650 284
rect -50 216 -45 250
rect 645 216 650 250
rect -50 182 -37 216
rect 637 182 650 216
rect -50 148 -45 182
rect 645 148 650 182
rect -50 114 -37 148
rect 637 114 650 148
rect -50 80 -45 114
rect 645 80 650 114
rect -50 46 -37 80
rect 637 46 650 80
rect -50 0 -45 46
rect 645 0 650 46
<< nwell >>
rect -81 -36 681 1386
<< pmos >>
rect 0 0 600 1350
<< pdiff >>
rect -45 1304 0 1350
rect -11 1270 0 1304
rect -45 1236 0 1270
rect -11 1202 0 1236
rect -45 1168 0 1202
rect -11 1134 0 1168
rect -45 1100 0 1134
rect -11 1066 0 1100
rect -45 1032 0 1066
rect -11 998 0 1032
rect -45 964 0 998
rect -11 930 0 964
rect -45 896 0 930
rect -11 862 0 896
rect -45 828 0 862
rect -11 794 0 828
rect -45 760 0 794
rect -11 726 0 760
rect -45 692 0 726
rect -11 658 0 692
rect -45 624 0 658
rect -11 590 0 624
rect -45 556 0 590
rect -11 522 0 556
rect -45 488 0 522
rect -11 454 0 488
rect -45 420 0 454
rect -11 386 0 420
rect -45 352 0 386
rect -11 318 0 352
rect -45 284 0 318
rect -11 250 0 284
rect -45 216 0 250
rect -11 182 0 216
rect -45 148 0 182
rect -11 114 0 148
rect -45 80 0 114
rect -11 46 0 80
rect -45 0 0 46
rect 600 1304 645 1350
rect 600 1270 611 1304
rect 600 1236 645 1270
rect 600 1202 611 1236
rect 600 1168 645 1202
rect 600 1134 611 1168
rect 600 1100 645 1134
rect 600 1066 611 1100
rect 600 1032 645 1066
rect 600 998 611 1032
rect 600 964 645 998
rect 600 930 611 964
rect 600 896 645 930
rect 600 862 611 896
rect 600 828 645 862
rect 600 794 611 828
rect 600 760 645 794
rect 600 726 611 760
rect 600 692 645 726
rect 600 658 611 692
rect 600 624 645 658
rect 600 590 611 624
rect 600 556 645 590
rect 600 522 611 556
rect 600 488 645 522
rect 600 454 611 488
rect 600 420 645 454
rect 600 386 611 420
rect 600 352 645 386
rect 600 318 611 352
rect 600 284 645 318
rect 600 250 611 284
rect 600 216 645 250
rect 600 182 611 216
rect 600 148 645 182
rect 600 114 611 148
rect 600 80 645 114
rect 600 46 611 80
rect 600 0 645 46
<< pdiffc >>
rect -45 1270 -11 1304
rect -45 1202 -11 1236
rect -45 1134 -11 1168
rect -45 1066 -11 1100
rect -45 998 -11 1032
rect -45 930 -11 964
rect -45 862 -11 896
rect -45 794 -11 828
rect -45 726 -11 760
rect -45 658 -11 692
rect -45 590 -11 624
rect -45 522 -11 556
rect -45 454 -11 488
rect -45 386 -11 420
rect -45 318 -11 352
rect -45 250 -11 284
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect 611 1270 645 1304
rect 611 1202 645 1236
rect 611 1134 645 1168
rect 611 1066 645 1100
rect 611 998 645 1032
rect 611 930 645 964
rect 611 862 645 896
rect 611 794 645 828
rect 611 726 645 760
rect 611 658 645 692
rect 611 590 645 624
rect 611 522 645 556
rect 611 454 645 488
rect 611 386 645 420
rect 611 318 645 352
rect 611 250 645 284
rect 611 182 645 216
rect 611 114 645 148
rect 611 46 645 80
<< poly >>
rect 0 1350 600 1380
rect 0 -48 600 0
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< polycont >>
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< locali >>
rect -45 1304 -11 1350
rect -45 1236 -11 1270
rect -45 1168 -11 1202
rect -45 1100 -11 1134
rect -45 1032 -11 1066
rect -45 964 -11 998
rect -45 896 -11 930
rect -45 828 -11 862
rect -45 760 -11 794
rect -45 692 -11 726
rect -45 624 -11 658
rect -45 556 -11 590
rect -45 488 -11 522
rect -45 420 -11 454
rect -45 352 -11 386
rect -45 284 -11 318
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 0 -11 46
rect 611 1304 645 1350
rect 611 1236 645 1270
rect 611 1168 645 1202
rect 611 1100 645 1134
rect 611 1032 645 1066
rect 611 964 645 998
rect 611 896 645 930
rect 611 828 645 862
rect 611 760 645 794
rect 611 692 645 726
rect 611 624 645 658
rect 611 556 645 590
rect 611 488 645 522
rect 611 420 645 454
rect 611 352 645 386
rect 611 284 645 318
rect 611 216 645 250
rect 611 148 645 182
rect 611 80 645 114
rect 611 0 645 46
rect 0 -48 600 -42
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -88 600 -82
<< viali >>
rect 16 -82 50 -48
rect 93 -82 127 -48
rect 170 -82 204 -48
rect 246 -82 280 -48
rect 322 -82 356 -48
rect 398 -82 432 -48
rect 474 -82 508 -48
rect 550 -82 584 -48
<< metal1 >>
rect 0 -48 600 -38
rect 0 -82 16 -48
rect 50 -82 93 -48
rect 127 -82 170 -48
rect 204 -82 246 -48
rect 280 -82 322 -48
rect 356 -82 398 -48
rect 432 -82 474 -48
rect 508 -82 550 -48
rect 584 -82 600 -48
rect 0 -92 600 -82
<< end >>
