magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 0 -21 200
<< pwell >>
rect -47 -154 109 226
<< nmos >>
rect 0 0 30 200
<< ndiff >>
rect -21 0 0 200
rect 30 151 83 200
rect 30 117 41 151
rect 75 117 83 151
rect 30 83 83 117
rect 30 49 41 83
rect 75 49 83 83
rect 30 0 83 49
<< ndiffc >>
rect 41 117 75 151
rect 41 49 75 83
<< psubdiff >>
rect -21 -82 83 -70
rect -21 -116 14 -82
rect 48 -116 83 -82
rect -21 -128 83 -116
<< psubdiffcont >>
rect 14 -116 48 -82
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect 41 151 75 200
rect 41 83 75 117
rect 41 0 75 49
rect -19 -82 81 -72
rect -19 -116 14 -82
rect 48 -116 81 -82
rect -19 -126 81 -116
<< viali >>
rect 14 -116 48 -82
<< metal1 >>
rect -19 -82 81 -72
rect -19 -116 14 -82
rect 48 -116 81 -82
rect -19 -126 81 -116
<< end >>
