magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -17 -17 17 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -37 17 37 23
rect -37 -17 -17 17
rect 17 -17 37 17
rect -37 -23 37 -17
<< end >>
