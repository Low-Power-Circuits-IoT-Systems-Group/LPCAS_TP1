magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -29 17 29 27
rect -29 -17 -17 17
rect -29 -27 29 -17
<< locali >>
rect -27 -17 -17 17
rect 17 -17 27 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -29 17 29 27
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -27 29 -17
<< end >>
