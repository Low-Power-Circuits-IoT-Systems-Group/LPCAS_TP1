magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 1969 -45 2000
rect -50 1935 -37 1969
rect -50 1901 -45 1935
rect -50 1867 -37 1901
rect -50 1833 -45 1867
rect -50 1799 -37 1833
rect -50 1765 -45 1799
rect -50 1731 -37 1765
rect -50 1697 -45 1731
rect -50 1663 -37 1697
rect -50 1629 -45 1663
rect -50 1595 -37 1629
rect -50 1561 -45 1595
rect -50 1527 -37 1561
rect -50 1493 -45 1527
rect -50 1459 -37 1493
rect -50 1425 -45 1459
rect -50 1391 -37 1425
rect -50 1357 -45 1391
rect -50 1323 -37 1357
rect -50 1289 -45 1323
rect -50 1255 -37 1289
rect -50 1221 -45 1255
rect -50 1187 -37 1221
rect -50 1153 -45 1187
rect -50 1119 -37 1153
rect -50 1085 -45 1119
rect -50 1051 -37 1085
rect -50 1017 -45 1051
rect -50 983 -37 1017
rect -50 949 -45 983
rect -50 915 -37 949
rect -50 881 -45 915
rect -50 847 -37 881
rect -50 813 -45 847
rect -50 779 -37 813
rect -50 745 -45 779
rect -50 711 -37 745
rect -50 677 -45 711
rect -50 643 -37 677
rect -50 609 -45 643
rect -50 575 -37 609
rect -50 541 -45 575
rect -50 507 -37 541
rect -50 473 -45 507
rect -50 439 -37 473
rect -50 405 -45 439
rect -50 371 -37 405
rect -50 337 -45 371
rect -50 303 -37 337
rect -50 269 -45 303
rect -50 235 -37 269
rect -50 201 -45 235
rect -50 167 -37 201
rect -50 133 -45 167
rect -50 99 -37 133
rect -50 65 -45 99
rect -50 31 -37 65
rect -50 0 -45 31
<< pwell >>
rect -71 -154 109 2026
<< nmos >>
rect 0 0 30 2000
<< ndiff >>
rect -45 1969 0 2000
rect -11 1935 0 1969
rect -45 1901 0 1935
rect -11 1867 0 1901
rect -45 1833 0 1867
rect -11 1799 0 1833
rect -45 1765 0 1799
rect -11 1731 0 1765
rect -45 1697 0 1731
rect -11 1663 0 1697
rect -45 1629 0 1663
rect -11 1595 0 1629
rect -45 1561 0 1595
rect -11 1527 0 1561
rect -45 1493 0 1527
rect -11 1459 0 1493
rect -45 1425 0 1459
rect -11 1391 0 1425
rect -45 1357 0 1391
rect -11 1323 0 1357
rect -45 1289 0 1323
rect -11 1255 0 1289
rect -45 1221 0 1255
rect -11 1187 0 1221
rect -45 1153 0 1187
rect -11 1119 0 1153
rect -45 1085 0 1119
rect -11 1051 0 1085
rect -45 1017 0 1051
rect -11 983 0 1017
rect -45 949 0 983
rect -11 915 0 949
rect -45 881 0 915
rect -11 847 0 881
rect -45 813 0 847
rect -11 779 0 813
rect -45 745 0 779
rect -11 711 0 745
rect -45 677 0 711
rect -11 643 0 677
rect -45 609 0 643
rect -11 575 0 609
rect -45 541 0 575
rect -11 507 0 541
rect -45 473 0 507
rect -11 439 0 473
rect -45 405 0 439
rect -11 371 0 405
rect -45 337 0 371
rect -11 303 0 337
rect -45 269 0 303
rect -11 235 0 269
rect -45 201 0 235
rect -11 167 0 201
rect -45 133 0 167
rect -11 99 0 133
rect -45 65 0 99
rect -11 31 0 65
rect -45 0 0 31
rect 30 1969 83 2000
rect 30 1935 41 1969
rect 75 1935 83 1969
rect 30 1901 83 1935
rect 30 1867 41 1901
rect 75 1867 83 1901
rect 30 1833 83 1867
rect 30 1799 41 1833
rect 75 1799 83 1833
rect 30 1765 83 1799
rect 30 1731 41 1765
rect 75 1731 83 1765
rect 30 1697 83 1731
rect 30 1663 41 1697
rect 75 1663 83 1697
rect 30 1629 83 1663
rect 30 1595 41 1629
rect 75 1595 83 1629
rect 30 1561 83 1595
rect 30 1527 41 1561
rect 75 1527 83 1561
rect 30 1493 83 1527
rect 30 1459 41 1493
rect 75 1459 83 1493
rect 30 1425 83 1459
rect 30 1391 41 1425
rect 75 1391 83 1425
rect 30 1357 83 1391
rect 30 1323 41 1357
rect 75 1323 83 1357
rect 30 1289 83 1323
rect 30 1255 41 1289
rect 75 1255 83 1289
rect 30 1221 83 1255
rect 30 1187 41 1221
rect 75 1187 83 1221
rect 30 1153 83 1187
rect 30 1119 41 1153
rect 75 1119 83 1153
rect 30 1085 83 1119
rect 30 1051 41 1085
rect 75 1051 83 1085
rect 30 1017 83 1051
rect 30 983 41 1017
rect 75 983 83 1017
rect 30 949 83 983
rect 30 915 41 949
rect 75 915 83 949
rect 30 881 83 915
rect 30 847 41 881
rect 75 847 83 881
rect 30 813 83 847
rect 30 779 41 813
rect 75 779 83 813
rect 30 745 83 779
rect 30 711 41 745
rect 75 711 83 745
rect 30 677 83 711
rect 30 643 41 677
rect 75 643 83 677
rect 30 609 83 643
rect 30 575 41 609
rect 75 575 83 609
rect 30 541 83 575
rect 30 507 41 541
rect 75 507 83 541
rect 30 473 83 507
rect 30 439 41 473
rect 75 439 83 473
rect 30 405 83 439
rect 30 371 41 405
rect 75 371 83 405
rect 30 337 83 371
rect 30 303 41 337
rect 75 303 83 337
rect 30 269 83 303
rect 30 235 41 269
rect 75 235 83 269
rect 30 201 83 235
rect 30 167 41 201
rect 75 167 83 201
rect 30 133 83 167
rect 30 99 41 133
rect 75 99 83 133
rect 30 65 83 99
rect 30 31 41 65
rect 75 31 83 65
rect 30 0 83 31
<< ndiffc >>
rect -45 1935 -11 1969
rect -45 1867 -11 1901
rect -45 1799 -11 1833
rect -45 1731 -11 1765
rect -45 1663 -11 1697
rect -45 1595 -11 1629
rect -45 1527 -11 1561
rect -45 1459 -11 1493
rect -45 1391 -11 1425
rect -45 1323 -11 1357
rect -45 1255 -11 1289
rect -45 1187 -11 1221
rect -45 1119 -11 1153
rect -45 1051 -11 1085
rect -45 983 -11 1017
rect -45 915 -11 949
rect -45 847 -11 881
rect -45 779 -11 813
rect -45 711 -11 745
rect -45 643 -11 677
rect -45 575 -11 609
rect -45 507 -11 541
rect -45 439 -11 473
rect -45 371 -11 405
rect -45 303 -11 337
rect -45 235 -11 269
rect -45 167 -11 201
rect -45 99 -11 133
rect -45 31 -11 65
rect 41 1935 75 1969
rect 41 1867 75 1901
rect 41 1799 75 1833
rect 41 1731 75 1765
rect 41 1663 75 1697
rect 41 1595 75 1629
rect 41 1527 75 1561
rect 41 1459 75 1493
rect 41 1391 75 1425
rect 41 1323 75 1357
rect 41 1255 75 1289
rect 41 1187 75 1221
rect 41 1119 75 1153
rect 41 1051 75 1085
rect 41 983 75 1017
rect 41 915 75 949
rect 41 847 75 881
rect 41 779 75 813
rect 41 711 75 745
rect 41 643 75 677
rect 41 575 75 609
rect 41 507 75 541
rect 41 439 75 473
rect 41 371 75 405
rect 41 303 75 337
rect 41 235 75 269
rect 41 167 75 201
rect 41 99 75 133
rect 41 31 75 65
<< psubdiff >>
rect -45 -82 83 -70
rect -45 -116 2 -82
rect 36 -116 83 -82
rect -45 -128 83 -116
<< psubdiffcont >>
rect 2 -116 36 -82
<< poly >>
rect 0 2000 30 2030
rect 0 -30 30 0
<< locali >>
rect -45 1969 -11 2000
rect -45 1901 -11 1935
rect -45 1833 -11 1867
rect -45 1765 -11 1799
rect -45 1697 -11 1731
rect -45 1629 -11 1663
rect -45 1561 -11 1595
rect -45 1493 -11 1527
rect -45 1425 -11 1459
rect -45 1357 -11 1391
rect -45 1289 -11 1323
rect -45 1221 -11 1255
rect -45 1153 -11 1187
rect -45 1085 -11 1119
rect -45 1017 -11 1051
rect -45 949 -11 983
rect -45 881 -11 915
rect -45 813 -11 847
rect -45 745 -11 779
rect -45 677 -11 711
rect -45 609 -11 643
rect -45 541 -11 575
rect -45 473 -11 507
rect -45 405 -11 439
rect -45 337 -11 371
rect -45 269 -11 303
rect -45 201 -11 235
rect -45 133 -11 167
rect -45 65 -11 99
rect -45 0 -11 31
rect 41 1969 75 2000
rect 41 1901 75 1935
rect 41 1833 75 1867
rect 41 1765 75 1799
rect 41 1697 75 1731
rect 41 1629 75 1663
rect 41 1561 75 1595
rect 41 1493 75 1527
rect 41 1425 75 1459
rect 41 1357 75 1391
rect 41 1289 75 1323
rect 41 1221 75 1255
rect 41 1153 75 1187
rect 41 1085 75 1119
rect 41 1017 75 1051
rect 41 949 75 983
rect 41 881 75 915
rect 41 813 75 847
rect 41 745 75 779
rect 41 677 75 711
rect 41 609 75 643
rect 41 541 75 575
rect 41 473 75 507
rect 41 405 75 439
rect 41 337 75 371
rect 41 269 75 303
rect 41 201 75 235
rect 41 133 75 167
rect 41 65 75 99
rect 41 0 75 31
rect -43 -82 81 -72
rect -43 -116 2 -82
rect 36 -116 81 -82
rect -43 -126 81 -116
<< viali >>
rect 2 -116 36 -82
<< metal1 >>
rect -43 -82 81 -72
rect -43 -116 2 -82
rect 36 -116 81 -82
rect -43 -126 81 -116
<< end >>
