magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 51 0 80 200
<< nwell >>
rect -89 -36 87 362
<< pmos >>
rect 0 0 30 200
<< pdiff >>
rect -53 151 0 200
rect -53 117 -45 151
rect -11 117 0 151
rect -53 83 0 117
rect -53 49 -45 83
rect -11 49 0 83
rect -53 0 0 49
rect 30 0 51 200
<< pdiffc >>
rect -45 117 -11 151
rect -45 49 -11 83
<< nsubdiff >>
rect -53 314 51 326
rect -53 280 -18 314
rect 16 280 51 314
rect -53 268 51 280
<< nsubdiffcont >>
rect -18 280 16 314
<< poly >>
rect 0 200 30 230
rect 0 -30 30 0
<< locali >>
rect -51 314 49 324
rect -51 280 -18 314
rect 16 280 49 314
rect -51 270 49 280
rect -45 151 -11 200
rect -45 83 -11 117
rect -45 0 -11 49
<< viali >>
rect -18 280 16 314
<< metal1 >>
rect -51 314 49 324
rect -51 280 -18 314
rect 16 280 49 314
rect -51 270 49 280
<< end >>
