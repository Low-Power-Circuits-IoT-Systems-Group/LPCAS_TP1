magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< locali >>
rect -17 89 17 105
rect -17 17 17 55
rect -17 -55 17 -17
rect -17 -105 17 -89
<< viali >>
rect -17 55 17 89
rect -17 -17 17 17
rect -17 -89 17 -55
<< metal1 >>
rect -23 89 23 101
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -101 23 -89
<< end >>
