magic
tech sky130A
timestamp 1741700111
<< metal1 >>
rect -96 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 96 13
<< via1 >>
rect -93 -13 -67 13
rect -61 -13 -35 13
rect -29 -13 -3 13
rect 3 -13 29 13
rect 35 -13 61 13
rect 67 -13 93 13
<< metal2 >>
rect -96 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 96 13
<< end >>
