magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 545 471 550 500
rect 537 437 550 471
rect 545 403 550 437
rect 537 369 550 403
rect 545 335 550 369
rect 537 301 550 335
rect 545 267 550 301
rect 537 233 550 267
rect 545 199 550 233
rect 537 165 550 199
rect 545 131 550 165
rect 537 97 550 131
rect 545 63 550 97
rect 537 29 550 63
rect 545 0 550 29
<< pwell >>
rect -79 -26 571 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -53 471 0 500
rect -53 437 -45 471
rect -11 437 0 471
rect -53 403 0 437
rect -53 369 -45 403
rect -11 369 0 403
rect -53 335 0 369
rect -53 301 -45 335
rect -11 301 0 335
rect -53 267 0 301
rect -53 233 -45 267
rect -11 233 0 267
rect -53 199 0 233
rect -53 165 -45 199
rect -11 165 0 199
rect -53 131 0 165
rect -53 97 -45 131
rect -11 97 0 131
rect -53 63 0 97
rect -53 29 -45 63
rect -11 29 0 63
rect -53 0 0 29
rect 500 471 545 500
rect 500 437 511 471
rect 500 403 545 437
rect 500 369 511 403
rect 500 335 545 369
rect 500 301 511 335
rect 500 267 545 301
rect 500 233 511 267
rect 500 199 545 233
rect 500 165 511 199
rect 500 131 545 165
rect 500 97 511 131
rect 500 63 545 97
rect 500 29 511 63
rect 500 0 545 29
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
rect 511 437 545 471
rect 511 369 545 403
rect 511 301 545 335
rect 511 233 545 267
rect 511 165 545 199
rect 511 97 545 131
rect 511 29 545 63
<< poly >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 500 500 548
rect 0 -30 500 0
<< polycont >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< locali >>
rect 0 582 500 588
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 542 500 548
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect 511 471 545 500
rect 511 403 545 437
rect 511 335 545 369
rect 511 267 545 301
rect 511 199 545 233
rect 511 131 545 165
rect 511 63 545 97
rect 511 0 545 29
<< viali >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< metal1 >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 538 500 548
<< end >>
