magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 311 0 330 1400
<< pwell >>
rect -79 -26 337 1554
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -53 1363 0 1400
rect -53 1329 -45 1363
rect -11 1329 0 1363
rect -53 1295 0 1329
rect -53 1261 -45 1295
rect -11 1261 0 1295
rect -53 1227 0 1261
rect -53 1193 -45 1227
rect -11 1193 0 1227
rect -53 1159 0 1193
rect -53 1125 -45 1159
rect -11 1125 0 1159
rect -53 1091 0 1125
rect -53 1057 -45 1091
rect -11 1057 0 1091
rect -53 1023 0 1057
rect -53 989 -45 1023
rect -11 989 0 1023
rect -53 955 0 989
rect -53 921 -45 955
rect -11 921 0 955
rect -53 887 0 921
rect -53 853 -45 887
rect -11 853 0 887
rect -53 819 0 853
rect -53 785 -45 819
rect -11 785 0 819
rect -53 751 0 785
rect -53 717 -45 751
rect -11 717 0 751
rect -53 683 0 717
rect -53 649 -45 683
rect -11 649 0 683
rect -53 615 0 649
rect -53 581 -45 615
rect -11 581 0 615
rect -53 547 0 581
rect -53 513 -45 547
rect -11 513 0 547
rect -53 479 0 513
rect -53 445 -45 479
rect -11 445 0 479
rect -53 411 0 445
rect -53 377 -45 411
rect -11 377 0 411
rect -53 343 0 377
rect -53 309 -45 343
rect -11 309 0 343
rect -53 275 0 309
rect -53 241 -45 275
rect -11 241 0 275
rect -53 207 0 241
rect -53 173 -45 207
rect -11 173 0 207
rect -53 139 0 173
rect -53 105 -45 139
rect -11 105 0 139
rect -53 71 0 105
rect -53 37 -45 71
rect -11 37 0 71
rect -53 0 0 37
rect 300 0 311 1400
<< ndiffc >>
rect -45 1329 -11 1363
rect -45 1261 -11 1295
rect -45 1193 -11 1227
rect -45 1125 -11 1159
rect -45 1057 -11 1091
rect -45 989 -11 1023
rect -45 921 -11 955
rect -45 853 -11 887
rect -45 785 -11 819
rect -45 717 -11 751
rect -45 649 -11 683
rect -45 581 -11 615
rect -45 513 -11 547
rect -45 445 -11 479
rect -45 377 -11 411
rect -45 309 -11 343
rect -45 241 -11 275
rect -45 173 -11 207
rect -45 105 -11 139
rect -45 37 -11 71
<< psubdiff >>
rect -53 1516 311 1528
rect -53 1482 -24 1516
rect 10 1482 44 1516
rect 78 1482 112 1516
rect 146 1482 180 1516
rect 214 1482 248 1516
rect 282 1482 311 1516
rect -53 1470 311 1482
<< psubdiffcont >>
rect -24 1482 10 1516
rect 44 1482 78 1516
rect 112 1482 146 1516
rect 180 1482 214 1516
rect 248 1482 282 1516
<< poly >>
rect 0 1400 300 1430
rect 0 -48 300 0
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< polycont >>
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< locali >>
rect -51 1516 309 1526
rect -51 1482 -32 1516
rect 10 1482 40 1516
rect 78 1482 112 1516
rect 146 1482 180 1516
rect 218 1482 248 1516
rect 290 1482 309 1516
rect -51 1472 309 1482
rect -45 1363 -11 1400
rect -45 1295 -11 1329
rect -45 1227 -11 1261
rect -45 1159 -11 1193
rect -45 1091 -11 1125
rect -45 1023 -11 1057
rect -45 955 -11 989
rect -45 887 -11 921
rect -45 819 -11 853
rect -45 751 -11 785
rect -45 683 -11 717
rect -45 615 -11 649
rect -45 547 -11 581
rect -45 479 -11 513
rect -45 411 -11 445
rect -45 343 -11 377
rect -45 275 -11 309
rect -45 207 -11 241
rect -45 139 -11 173
rect -45 71 -11 105
rect -45 0 -11 37
rect 0 -48 300 -42
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -88 300 -82
<< viali >>
rect -32 1482 -24 1516
rect -24 1482 2 1516
rect 40 1482 44 1516
rect 44 1482 74 1516
rect 112 1482 146 1516
rect 184 1482 214 1516
rect 214 1482 218 1516
rect 256 1482 282 1516
rect 282 1482 290 1516
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< metal1 >>
rect -51 1516 309 1526
rect -51 1482 -32 1516
rect 2 1482 40 1516
rect 74 1482 112 1516
rect 146 1482 184 1516
rect 218 1482 256 1516
rect 290 1482 309 1516
rect -51 1472 309 1482
rect 0 -48 300 -38
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< end >>
