magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 471 -45 500
rect -50 437 -37 471
rect -50 403 -45 437
rect -50 369 -37 403
rect -50 335 -45 369
rect -50 301 -37 335
rect -50 267 -45 301
rect -50 233 -37 267
rect -50 199 -45 233
rect -50 165 -37 199
rect -50 131 -45 165
rect -50 97 -37 131
rect -50 63 -45 97
rect -50 29 -37 63
rect -50 0 -45 29
rect 511 0 550 500
<< pwell >>
rect -71 -154 537 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -45 471 0 500
rect -11 437 0 471
rect -45 403 0 437
rect -11 369 0 403
rect -45 335 0 369
rect -11 301 0 335
rect -45 267 0 301
rect -11 233 0 267
rect -45 199 0 233
rect -11 165 0 199
rect -45 131 0 165
rect -11 97 0 131
rect -45 63 0 97
rect -11 29 0 63
rect -45 0 0 29
rect 500 0 511 500
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
<< psubdiff >>
rect -45 -82 511 -70
rect -45 -116 12 -82
rect 46 -116 80 -82
rect 114 -116 148 -82
rect 182 -116 216 -82
rect 250 -116 284 -82
rect 318 -116 352 -82
rect 386 -116 420 -82
rect 454 -116 511 -82
rect -45 -128 511 -116
<< psubdiffcont >>
rect 12 -116 46 -82
rect 80 -116 114 -82
rect 148 -116 182 -82
rect 216 -116 250 -82
rect 284 -116 318 -82
rect 352 -116 386 -82
rect 420 -116 454 -82
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect -43 -82 509 -72
rect -43 -116 0 -82
rect 46 -116 72 -82
rect 114 -116 144 -82
rect 182 -116 216 -82
rect 250 -116 284 -82
rect 322 -116 352 -82
rect 394 -116 420 -82
rect 466 -116 509 -82
rect -43 -126 509 -116
<< viali >>
rect 0 -116 12 -82
rect 12 -116 34 -82
rect 72 -116 80 -82
rect 80 -116 106 -82
rect 144 -116 148 -82
rect 148 -116 178 -82
rect 216 -116 250 -82
rect 288 -116 318 -82
rect 318 -116 322 -82
rect 360 -116 386 -82
rect 386 -116 394 -82
rect 432 -116 454 -82
rect 454 -116 466 -82
<< metal1 >>
rect -43 -82 509 -72
rect -43 -116 0 -82
rect 34 -116 72 -82
rect 106 -116 144 -82
rect 178 -116 216 -82
rect 250 -116 288 -82
rect 322 -116 360 -82
rect 394 -116 432 -82
rect 466 -116 509 -82
rect -43 -126 509 -116
<< end >>
