magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -43 26 9 32
rect -43 -32 9 -26
<< via1 >>
rect -43 -26 9 26
<< metal2 >>
rect -45 26 11 37
rect -45 -26 -43 26
rect 9 -26 11 26
rect -45 -37 11 -26
<< end >>
