magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 511 0 550 500
<< pwell >>
rect -79 -154 537 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -53 471 0 500
rect -53 437 -45 471
rect -11 437 0 471
rect -53 403 0 437
rect -53 369 -45 403
rect -11 369 0 403
rect -53 335 0 369
rect -53 301 -45 335
rect -11 301 0 335
rect -53 267 0 301
rect -53 233 -45 267
rect -11 233 0 267
rect -53 199 0 233
rect -53 165 -45 199
rect -11 165 0 199
rect -53 131 0 165
rect -53 97 -45 131
rect -11 97 0 131
rect -53 63 0 97
rect -53 29 -45 63
rect -11 29 0 63
rect -53 0 0 29
rect 500 0 511 500
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
<< psubdiff >>
rect -53 -82 511 -70
rect -53 -116 -26 -82
rect 8 -116 42 -82
rect 76 -116 110 -82
rect 144 -116 178 -82
rect 212 -116 246 -82
rect 280 -116 314 -82
rect 348 -116 382 -82
rect 416 -116 450 -82
rect 484 -116 511 -82
rect -53 -128 511 -116
<< psubdiffcont >>
rect -26 -116 8 -82
rect 42 -116 76 -82
rect 110 -116 144 -82
rect 178 -116 212 -82
rect 246 -116 280 -82
rect 314 -116 348 -82
rect 382 -116 416 -82
rect 450 -116 484 -82
<< poly >>
rect 0 500 500 530
rect 0 -30 500 0
<< locali >>
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
rect -51 -82 509 -72
rect -51 -116 -26 -82
rect 30 -116 42 -82
rect 102 -116 110 -82
rect 174 -116 178 -82
rect 280 -116 284 -82
rect 348 -116 356 -82
rect 416 -116 428 -82
rect 484 -116 509 -82
rect -51 -126 509 -116
<< viali >>
rect -4 -116 8 -82
rect 8 -116 30 -82
rect 68 -116 76 -82
rect 76 -116 102 -82
rect 140 -116 144 -82
rect 144 -116 174 -82
rect 212 -116 246 -82
rect 284 -116 314 -82
rect 314 -116 318 -82
rect 356 -116 382 -82
rect 382 -116 390 -82
rect 428 -116 450 -82
rect 450 -116 462 -82
<< metal1 >>
rect -51 -82 509 -72
rect -51 -116 -4 -82
rect 30 -116 68 -82
rect 102 -116 140 -82
rect 174 -116 212 -82
rect 246 -116 284 -82
rect 318 -116 356 -82
rect 390 -116 428 -82
rect 462 -116 509 -82
rect -51 -126 509 -116
<< end >>
