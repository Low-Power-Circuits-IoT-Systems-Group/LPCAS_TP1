magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< metal1 >>
rect -101 -90 -90 90
rect 90 -90 101 90
<< via1 >>
rect -90 -90 90 90
<< metal2 >>
rect -101 -90 -90 90
rect 90 -90 101 90
<< end >>
