magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 41 0 80 2000
<< pwell >>
rect -79 -154 67 2026
<< nmos >>
rect 0 0 30 2000
<< ndiff >>
rect -53 1969 0 2000
rect -53 1935 -45 1969
rect -11 1935 0 1969
rect -53 1901 0 1935
rect -53 1867 -45 1901
rect -11 1867 0 1901
rect -53 1833 0 1867
rect -53 1799 -45 1833
rect -11 1799 0 1833
rect -53 1765 0 1799
rect -53 1731 -45 1765
rect -11 1731 0 1765
rect -53 1697 0 1731
rect -53 1663 -45 1697
rect -11 1663 0 1697
rect -53 1629 0 1663
rect -53 1595 -45 1629
rect -11 1595 0 1629
rect -53 1561 0 1595
rect -53 1527 -45 1561
rect -11 1527 0 1561
rect -53 1493 0 1527
rect -53 1459 -45 1493
rect -11 1459 0 1493
rect -53 1425 0 1459
rect -53 1391 -45 1425
rect -11 1391 0 1425
rect -53 1357 0 1391
rect -53 1323 -45 1357
rect -11 1323 0 1357
rect -53 1289 0 1323
rect -53 1255 -45 1289
rect -11 1255 0 1289
rect -53 1221 0 1255
rect -53 1187 -45 1221
rect -11 1187 0 1221
rect -53 1153 0 1187
rect -53 1119 -45 1153
rect -11 1119 0 1153
rect -53 1085 0 1119
rect -53 1051 -45 1085
rect -11 1051 0 1085
rect -53 1017 0 1051
rect -53 983 -45 1017
rect -11 983 0 1017
rect -53 949 0 983
rect -53 915 -45 949
rect -11 915 0 949
rect -53 881 0 915
rect -53 847 -45 881
rect -11 847 0 881
rect -53 813 0 847
rect -53 779 -45 813
rect -11 779 0 813
rect -53 745 0 779
rect -53 711 -45 745
rect -11 711 0 745
rect -53 677 0 711
rect -53 643 -45 677
rect -11 643 0 677
rect -53 609 0 643
rect -53 575 -45 609
rect -11 575 0 609
rect -53 541 0 575
rect -53 507 -45 541
rect -11 507 0 541
rect -53 473 0 507
rect -53 439 -45 473
rect -11 439 0 473
rect -53 405 0 439
rect -53 371 -45 405
rect -11 371 0 405
rect -53 337 0 371
rect -53 303 -45 337
rect -11 303 0 337
rect -53 269 0 303
rect -53 235 -45 269
rect -11 235 0 269
rect -53 201 0 235
rect -53 167 -45 201
rect -11 167 0 201
rect -53 133 0 167
rect -53 99 -45 133
rect -11 99 0 133
rect -53 65 0 99
rect -53 31 -45 65
rect -11 31 0 65
rect -53 0 0 31
rect 30 0 41 2000
<< ndiffc >>
rect -45 1935 -11 1969
rect -45 1867 -11 1901
rect -45 1799 -11 1833
rect -45 1731 -11 1765
rect -45 1663 -11 1697
rect -45 1595 -11 1629
rect -45 1527 -11 1561
rect -45 1459 -11 1493
rect -45 1391 -11 1425
rect -45 1323 -11 1357
rect -45 1255 -11 1289
rect -45 1187 -11 1221
rect -45 1119 -11 1153
rect -45 1051 -11 1085
rect -45 983 -11 1017
rect -45 915 -11 949
rect -45 847 -11 881
rect -45 779 -11 813
rect -45 711 -11 745
rect -45 643 -11 677
rect -45 575 -11 609
rect -45 507 -11 541
rect -45 439 -11 473
rect -45 371 -11 405
rect -45 303 -11 337
rect -45 235 -11 269
rect -45 167 -11 201
rect -45 99 -11 133
rect -45 31 -11 65
<< psubdiff >>
rect -53 -82 41 -70
rect -53 -116 -23 -82
rect 11 -116 41 -82
rect -53 -128 41 -116
<< psubdiffcont >>
rect -23 -116 11 -82
<< poly >>
rect 0 2000 30 2030
rect 0 -30 30 0
<< locali >>
rect -45 1969 -11 2000
rect -45 1901 -11 1935
rect -45 1833 -11 1867
rect -45 1765 -11 1799
rect -45 1697 -11 1731
rect -45 1629 -11 1663
rect -45 1561 -11 1595
rect -45 1493 -11 1527
rect -45 1425 -11 1459
rect -45 1357 -11 1391
rect -45 1289 -11 1323
rect -45 1221 -11 1255
rect -45 1153 -11 1187
rect -45 1085 -11 1119
rect -45 1017 -11 1051
rect -45 949 -11 983
rect -45 881 -11 915
rect -45 813 -11 847
rect -45 745 -11 779
rect -45 677 -11 711
rect -45 609 -11 643
rect -45 541 -11 575
rect -45 473 -11 507
rect -45 405 -11 439
rect -45 337 -11 371
rect -45 269 -11 303
rect -45 201 -11 235
rect -45 133 -11 167
rect -45 65 -11 99
rect -45 0 -11 31
rect -51 -82 39 -72
rect -51 -116 -23 -82
rect 11 -116 39 -82
rect -51 -126 39 -116
<< viali >>
rect -23 -116 11 -82
<< metal1 >>
rect -51 -82 39 -72
rect -51 -116 -23 -82
rect 11 -116 39 -82
rect -51 -126 39 -116
<< end >>
