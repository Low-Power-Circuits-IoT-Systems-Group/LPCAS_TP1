magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< nwell >>
rect -236 -36 1089 146
<< pmos >>
rect 0 0 1000 110
<< pdiff >>
rect -53 72 0 110
rect -53 38 -45 72
rect -11 38 0 72
rect -53 0 0 38
rect 1000 72 1053 110
rect 1000 38 1011 72
rect 1045 38 1053 72
rect 1000 0 1053 38
<< pdiffc >>
rect -45 38 -11 72
rect 1011 38 1045 72
<< nsubdiff >>
rect -200 72 -107 110
rect -200 38 -171 72
rect -137 38 -107 72
rect -200 0 -107 38
<< nsubdiffcont >>
rect -171 38 -137 72
<< poly >>
rect 0 110 1000 140
rect 0 -48 1000 0
rect 0 -82 16 -48
rect 50 -82 88 -48
rect 122 -82 160 -48
rect 194 -82 232 -48
rect 266 -82 304 -48
rect 338 -82 376 -48
rect 410 -82 448 -48
rect 482 -82 520 -48
rect 554 -82 592 -48
rect 626 -82 664 -48
rect 698 -82 736 -48
rect 770 -82 808 -48
rect 842 -82 879 -48
rect 913 -82 950 -48
rect 984 -82 1000 -48
rect 0 -92 1000 -82
<< polycont >>
rect 16 -82 50 -48
rect 88 -82 122 -48
rect 160 -82 194 -48
rect 232 -82 266 -48
rect 304 -82 338 -48
rect 376 -82 410 -48
rect 448 -82 482 -48
rect 520 -82 554 -48
rect 592 -82 626 -48
rect 664 -82 698 -48
rect 736 -82 770 -48
rect 808 -82 842 -48
rect 879 -82 913 -48
rect 950 -82 984 -48
<< locali >>
rect -198 72 -109 110
rect -198 38 -171 72
rect -137 38 -109 72
rect -198 0 -109 38
rect -45 72 -11 110
rect -45 0 -11 38
rect 1011 72 1045 110
rect 1011 0 1045 38
rect 0 -48 1000 -42
rect 0 -82 16 -48
rect 50 -82 88 -48
rect 128 -82 160 -48
rect 206 -82 232 -48
rect 284 -82 304 -48
rect 362 -82 376 -48
rect 440 -82 448 -48
rect 482 -82 484 -48
rect 518 -82 520 -48
rect 554 -82 562 -48
rect 626 -82 640 -48
rect 698 -82 718 -48
rect 770 -82 796 -48
rect 842 -82 873 -48
rect 913 -82 950 -48
rect 984 -82 1000 -48
rect 0 -88 1000 -82
<< viali >>
rect -171 38 -137 72
rect 16 -82 50 -48
rect 94 -82 122 -48
rect 122 -82 128 -48
rect 172 -82 194 -48
rect 194 -82 206 -48
rect 250 -82 266 -48
rect 266 -82 284 -48
rect 328 -82 338 -48
rect 338 -82 362 -48
rect 406 -82 410 -48
rect 410 -82 440 -48
rect 484 -82 518 -48
rect 562 -82 592 -48
rect 592 -82 596 -48
rect 640 -82 664 -48
rect 664 -82 674 -48
rect 718 -82 736 -48
rect 736 -82 752 -48
rect 796 -82 808 -48
rect 808 -82 830 -48
rect 873 -82 879 -48
rect 879 -82 907 -48
rect 950 -82 984 -48
<< metal1 >>
rect -198 72 -109 110
rect -198 38 -171 72
rect -137 38 -109 72
rect -198 0 -109 38
rect 0 -48 1000 -38
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 328 -48
rect 362 -82 406 -48
rect 440 -82 484 -48
rect 518 -82 562 -48
rect 596 -82 640 -48
rect 674 -82 718 -48
rect 752 -82 796 -48
rect 830 -82 873 -48
rect 907 -82 950 -48
rect 984 -82 1000 -48
rect 0 -92 1000 -82
<< end >>
