magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 1969 -45 2000
rect -50 1935 -37 1969
rect -50 1901 -45 1935
rect -50 1867 -37 1901
rect -50 1833 -45 1867
rect -50 1799 -37 1833
rect -50 1765 -45 1799
rect -50 1731 -37 1765
rect -50 1697 -45 1731
rect -50 1663 -37 1697
rect -50 1629 -45 1663
rect -50 1595 -37 1629
rect -50 1561 -45 1595
rect -50 1527 -37 1561
rect -50 1493 -45 1527
rect -50 1459 -37 1493
rect -50 1425 -45 1459
rect -50 1391 -37 1425
rect -50 1357 -45 1391
rect -50 1323 -37 1357
rect -50 1289 -45 1323
rect -50 1255 -37 1289
rect -50 1221 -45 1255
rect -50 1187 -37 1221
rect -50 1153 -45 1187
rect -50 1119 -37 1153
rect -50 1085 -45 1119
rect -50 1051 -37 1085
rect -50 1017 -45 1051
rect -50 983 -37 1017
rect -50 949 -45 983
rect -50 915 -37 949
rect -50 881 -45 915
rect -50 847 -37 881
rect -50 813 -45 847
rect -50 779 -37 813
rect -50 745 -45 779
rect -50 711 -37 745
rect -50 677 -45 711
rect -50 643 -37 677
rect -50 609 -45 643
rect -50 575 -37 609
rect -50 541 -45 575
rect -50 507 -37 541
rect -50 473 -45 507
rect -50 439 -37 473
rect -50 405 -45 439
rect -50 371 -37 405
rect -50 337 -45 371
rect -50 303 -37 337
rect -50 269 -45 303
rect -50 235 -37 269
rect -50 201 -45 235
rect -50 167 -37 201
rect -50 133 -45 167
rect -50 99 -37 133
rect -50 65 -45 99
rect -50 31 -37 65
rect -50 0 -45 31
rect 41 0 80 2000
<< pwell >>
rect -71 -154 67 2026
<< nmos >>
rect 0 0 30 2000
<< ndiff >>
rect -45 1969 0 2000
rect -11 1935 0 1969
rect -45 1901 0 1935
rect -11 1867 0 1901
rect -45 1833 0 1867
rect -11 1799 0 1833
rect -45 1765 0 1799
rect -11 1731 0 1765
rect -45 1697 0 1731
rect -11 1663 0 1697
rect -45 1629 0 1663
rect -11 1595 0 1629
rect -45 1561 0 1595
rect -11 1527 0 1561
rect -45 1493 0 1527
rect -11 1459 0 1493
rect -45 1425 0 1459
rect -11 1391 0 1425
rect -45 1357 0 1391
rect -11 1323 0 1357
rect -45 1289 0 1323
rect -11 1255 0 1289
rect -45 1221 0 1255
rect -11 1187 0 1221
rect -45 1153 0 1187
rect -11 1119 0 1153
rect -45 1085 0 1119
rect -11 1051 0 1085
rect -45 1017 0 1051
rect -11 983 0 1017
rect -45 949 0 983
rect -11 915 0 949
rect -45 881 0 915
rect -11 847 0 881
rect -45 813 0 847
rect -11 779 0 813
rect -45 745 0 779
rect -11 711 0 745
rect -45 677 0 711
rect -11 643 0 677
rect -45 609 0 643
rect -11 575 0 609
rect -45 541 0 575
rect -11 507 0 541
rect -45 473 0 507
rect -11 439 0 473
rect -45 405 0 439
rect -11 371 0 405
rect -45 337 0 371
rect -11 303 0 337
rect -45 269 0 303
rect -11 235 0 269
rect -45 201 0 235
rect -11 167 0 201
rect -45 133 0 167
rect -11 99 0 133
rect -45 65 0 99
rect -11 31 0 65
rect -45 0 0 31
rect 30 0 41 2000
<< ndiffc >>
rect -45 1935 -11 1969
rect -45 1867 -11 1901
rect -45 1799 -11 1833
rect -45 1731 -11 1765
rect -45 1663 -11 1697
rect -45 1595 -11 1629
rect -45 1527 -11 1561
rect -45 1459 -11 1493
rect -45 1391 -11 1425
rect -45 1323 -11 1357
rect -45 1255 -11 1289
rect -45 1187 -11 1221
rect -45 1119 -11 1153
rect -45 1051 -11 1085
rect -45 983 -11 1017
rect -45 915 -11 949
rect -45 847 -11 881
rect -45 779 -11 813
rect -45 711 -11 745
rect -45 643 -11 677
rect -45 575 -11 609
rect -45 507 -11 541
rect -45 439 -11 473
rect -45 371 -11 405
rect -45 303 -11 337
rect -45 235 -11 269
rect -45 167 -11 201
rect -45 99 -11 133
rect -45 31 -11 65
<< psubdiff >>
rect -45 -82 41 -70
rect -45 -116 -19 -82
rect 15 -116 41 -82
rect -45 -128 41 -116
<< psubdiffcont >>
rect -19 -116 15 -82
<< poly >>
rect 0 2000 30 2030
rect 0 -30 30 0
<< locali >>
rect -45 1969 -11 2000
rect -45 1901 -11 1935
rect -45 1833 -11 1867
rect -45 1765 -11 1799
rect -45 1697 -11 1731
rect -45 1629 -11 1663
rect -45 1561 -11 1595
rect -45 1493 -11 1527
rect -45 1425 -11 1459
rect -45 1357 -11 1391
rect -45 1289 -11 1323
rect -45 1221 -11 1255
rect -45 1153 -11 1187
rect -45 1085 -11 1119
rect -45 1017 -11 1051
rect -45 949 -11 983
rect -45 881 -11 915
rect -45 813 -11 847
rect -45 745 -11 779
rect -45 677 -11 711
rect -45 609 -11 643
rect -45 541 -11 575
rect -45 473 -11 507
rect -45 405 -11 439
rect -45 337 -11 371
rect -45 269 -11 303
rect -45 201 -11 235
rect -45 133 -11 167
rect -45 65 -11 99
rect -45 0 -11 31
rect -43 -82 39 -72
rect -43 -116 -19 -82
rect 15 -116 39 -82
rect -43 -126 39 -116
<< viali >>
rect -19 -116 15 -82
<< metal1 >>
rect -43 -82 39 -72
rect -43 -116 -19 -82
rect 15 -116 39 -82
rect -43 -126 39 -116
<< end >>
