magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< locali >>
rect -17 -19 17 19
<< viali >>
rect -17 19 17 53
rect -17 -53 17 -19
<< metal1 >>
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
<< end >>
