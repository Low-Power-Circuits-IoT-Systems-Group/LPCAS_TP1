magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 471 -45 500
rect -50 437 -37 471
rect -50 403 -45 437
rect -50 369 -37 403
rect -50 335 -45 369
rect -50 301 -37 335
rect -50 267 -45 301
rect -50 233 -37 267
rect -50 199 -45 233
rect -50 165 -37 199
rect -50 131 -45 165
rect -50 97 -37 131
rect -50 63 -45 97
rect -50 29 -37 63
rect -50 0 -45 29
rect 511 0 550 500
<< pwell >>
rect -71 -26 537 526
<< nmos >>
rect 0 0 500 500
<< ndiff >>
rect -45 471 0 500
rect -11 437 0 471
rect -45 403 0 437
rect -11 369 0 403
rect -45 335 0 369
rect -11 301 0 335
rect -45 267 0 301
rect -11 233 0 267
rect -45 199 0 233
rect -11 165 0 199
rect -45 131 0 165
rect -11 97 0 131
rect -45 63 0 97
rect -11 29 0 63
rect -45 0 0 29
rect 500 0 511 500
<< ndiffc >>
rect -45 437 -11 471
rect -45 369 -11 403
rect -45 301 -11 335
rect -45 233 -11 267
rect -45 165 -11 199
rect -45 97 -11 131
rect -45 29 -11 63
<< poly >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 500 500 548
rect 0 -30 500 0
<< polycont >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< locali >>
rect 0 582 500 588
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 542 500 548
rect -45 471 -11 500
rect -45 403 -11 437
rect -45 335 -11 369
rect -45 267 -11 301
rect -45 199 -11 233
rect -45 131 -11 165
rect -45 63 -11 97
rect -45 0 -11 29
<< viali >>
rect 16 548 50 582
rect 89 548 123 582
rect 162 548 196 582
rect 234 548 268 582
rect 306 548 340 582
rect 378 548 412 582
rect 450 548 484 582
<< metal1 >>
rect 0 582 500 592
rect 0 548 16 582
rect 50 548 89 582
rect 123 548 162 582
rect 196 548 234 582
rect 268 548 306 582
rect 340 548 378 582
rect 412 548 450 582
rect 484 548 500 582
rect 0 538 500 548
<< end >>
