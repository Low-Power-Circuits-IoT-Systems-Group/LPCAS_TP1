magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect 337 1329 345 1363
rect 337 1261 345 1295
rect 337 1193 345 1227
rect 337 1125 345 1159
rect 337 1057 345 1091
rect 337 989 345 1023
rect 337 921 345 955
rect 337 853 345 887
rect 337 785 345 819
rect 337 717 345 751
rect 337 649 345 683
rect 337 581 345 615
rect 337 513 345 547
rect 337 445 345 479
rect 337 377 345 411
rect 337 309 345 343
rect 337 241 345 275
rect 337 173 345 207
rect 337 105 345 139
rect 337 37 345 71
<< pwell >>
rect -79 -26 371 1554
<< nmoslvt >>
rect 0 0 300 1400
<< ndiff >>
rect -53 1363 0 1400
rect -53 1329 -45 1363
rect -11 1329 0 1363
rect -53 1295 0 1329
rect -53 1261 -45 1295
rect -11 1261 0 1295
rect -53 1227 0 1261
rect -53 1193 -45 1227
rect -11 1193 0 1227
rect -53 1159 0 1193
rect -53 1125 -45 1159
rect -11 1125 0 1159
rect -53 1091 0 1125
rect -53 1057 -45 1091
rect -11 1057 0 1091
rect -53 1023 0 1057
rect -53 989 -45 1023
rect -11 989 0 1023
rect -53 955 0 989
rect -53 921 -45 955
rect -11 921 0 955
rect -53 887 0 921
rect -53 853 -45 887
rect -11 853 0 887
rect -53 819 0 853
rect -53 785 -45 819
rect -11 785 0 819
rect -53 751 0 785
rect -53 717 -45 751
rect -11 717 0 751
rect -53 683 0 717
rect -53 649 -45 683
rect -11 649 0 683
rect -53 615 0 649
rect -53 581 -45 615
rect -11 581 0 615
rect -53 547 0 581
rect -53 513 -45 547
rect -11 513 0 547
rect -53 479 0 513
rect -53 445 -45 479
rect -11 445 0 479
rect -53 411 0 445
rect -53 377 -45 411
rect -11 377 0 411
rect -53 343 0 377
rect -53 309 -45 343
rect -11 309 0 343
rect -53 275 0 309
rect -53 241 -45 275
rect -11 241 0 275
rect -53 207 0 241
rect -53 173 -45 207
rect -11 173 0 207
rect -53 139 0 173
rect -53 105 -45 139
rect -11 105 0 139
rect -53 71 0 105
rect -53 37 -45 71
rect -11 37 0 71
rect -53 0 0 37
rect 300 1363 345 1400
rect 300 1329 311 1363
rect 300 1295 345 1329
rect 300 1261 311 1295
rect 300 1227 345 1261
rect 300 1193 311 1227
rect 300 1159 345 1193
rect 300 1125 311 1159
rect 300 1091 345 1125
rect 300 1057 311 1091
rect 300 1023 345 1057
rect 300 989 311 1023
rect 300 955 345 989
rect 300 921 311 955
rect 300 887 345 921
rect 300 853 311 887
rect 300 819 345 853
rect 300 785 311 819
rect 300 751 345 785
rect 300 717 311 751
rect 300 683 345 717
rect 300 649 311 683
rect 300 615 345 649
rect 300 581 311 615
rect 300 547 345 581
rect 300 513 311 547
rect 300 479 345 513
rect 300 445 311 479
rect 300 411 345 445
rect 300 377 311 411
rect 300 343 345 377
rect 300 309 311 343
rect 300 275 345 309
rect 300 241 311 275
rect 300 207 345 241
rect 300 173 311 207
rect 300 139 345 173
rect 300 105 311 139
rect 300 71 345 105
rect 300 37 311 71
rect 300 0 345 37
<< ndiffc >>
rect -45 1329 -11 1363
rect -45 1261 -11 1295
rect -45 1193 -11 1227
rect -45 1125 -11 1159
rect -45 1057 -11 1091
rect -45 989 -11 1023
rect -45 921 -11 955
rect -45 853 -11 887
rect -45 785 -11 819
rect -45 717 -11 751
rect -45 649 -11 683
rect -45 581 -11 615
rect -45 513 -11 547
rect -45 445 -11 479
rect -45 377 -11 411
rect -45 309 -11 343
rect -45 241 -11 275
rect -45 173 -11 207
rect -45 105 -11 139
rect -45 37 -11 71
rect 311 1329 345 1363
rect 311 1261 345 1295
rect 311 1193 345 1227
rect 311 1125 345 1159
rect 311 1057 345 1091
rect 311 989 345 1023
rect 311 921 345 955
rect 311 853 345 887
rect 311 785 345 819
rect 311 717 345 751
rect 311 649 345 683
rect 311 581 345 615
rect 311 513 345 547
rect 311 445 345 479
rect 311 377 345 411
rect 311 309 345 343
rect 311 241 345 275
rect 311 173 345 207
rect 311 105 345 139
rect 311 37 345 71
<< psubdiff >>
rect -53 1516 345 1528
rect -53 1482 -7 1516
rect 27 1482 61 1516
rect 95 1482 129 1516
rect 163 1482 197 1516
rect 231 1482 265 1516
rect 299 1482 345 1516
rect -53 1470 345 1482
<< psubdiffcont >>
rect -7 1482 27 1516
rect 61 1482 95 1516
rect 129 1482 163 1516
rect 197 1482 231 1516
rect 265 1482 299 1516
<< poly >>
rect 0 1400 300 1430
rect 0 -48 300 0
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< polycont >>
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< locali >>
rect -51 1516 343 1526
rect -51 1482 -15 1516
rect 27 1482 57 1516
rect 95 1482 129 1516
rect 163 1482 197 1516
rect 235 1482 265 1516
rect 307 1482 343 1516
rect -51 1472 343 1482
rect -45 1363 -11 1400
rect -45 1295 -11 1329
rect -45 1227 -11 1261
rect -45 1159 -11 1193
rect -45 1091 -11 1125
rect -45 1023 -11 1057
rect -45 955 -11 989
rect -45 887 -11 921
rect -45 819 -11 853
rect -45 751 -11 785
rect -45 683 -11 717
rect -45 615 -11 649
rect -45 547 -11 581
rect -45 479 -11 513
rect -45 411 -11 445
rect -45 343 -11 377
rect -45 275 -11 309
rect -45 207 -11 241
rect -45 139 -11 173
rect -45 71 -11 105
rect -45 0 -11 37
rect 311 1363 345 1400
rect 311 1295 345 1329
rect 311 1227 345 1261
rect 311 1159 345 1193
rect 311 1091 345 1125
rect 311 1023 345 1057
rect 311 955 345 989
rect 311 887 345 921
rect 311 819 345 853
rect 311 751 345 785
rect 311 683 345 717
rect 311 615 345 649
rect 311 547 345 581
rect 311 479 345 513
rect 311 411 345 445
rect 311 343 345 377
rect 311 275 345 309
rect 311 207 345 241
rect 311 139 345 173
rect 311 71 345 105
rect 311 0 345 37
rect 0 -48 300 -42
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -88 300 -82
<< viali >>
rect -15 1482 -7 1516
rect -7 1482 19 1516
rect 57 1482 61 1516
rect 61 1482 91 1516
rect 129 1482 163 1516
rect 201 1482 231 1516
rect 231 1482 235 1516
rect 273 1482 299 1516
rect 299 1482 307 1516
rect 16 -82 50 -48
rect 94 -82 128 -48
rect 172 -82 206 -48
rect 250 -82 284 -48
<< metal1 >>
rect -51 1516 343 1526
rect -51 1482 -15 1516
rect 19 1482 57 1516
rect 91 1482 129 1516
rect 163 1482 201 1516
rect 235 1482 273 1516
rect 307 1482 343 1516
rect -51 1472 343 1482
rect 0 -48 300 -38
rect 0 -82 16 -48
rect 50 -82 94 -48
rect 128 -82 172 -48
rect 206 -82 250 -48
rect 284 -82 300 -48
rect 0 -92 300 -82
<< end >>
