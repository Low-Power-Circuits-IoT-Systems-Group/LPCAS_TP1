magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< error_p >>
rect -50 28 16 33
rect -50 -28 -45 28
rect -50 -33 16 -28
<< metal2 >>
rect -45 28 11 37
rect -45 -37 11 -28
<< via2 >>
rect -45 -28 11 28
<< metal3 >>
rect -50 28 16 33
rect -50 -28 -45 28
rect 11 -28 16 28
rect -50 -33 16 -28
<< end >>
