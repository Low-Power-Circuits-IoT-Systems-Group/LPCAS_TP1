VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_LPCAS_TP1
  CLASS BLOCK ;
  FOREIGN tt_um_LPCAS_TP1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 18.150000 ;
    ANTENNADIFFAREA 15.650000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNADIFFAREA 7.542800 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNAGATEAREA 32.250000 ;
    ANTENNADIFFAREA 117.460548 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 7.500000 ;
    ANTENNADIFFAREA 10.934999 ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 2.950000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.200 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    ANTENNADIFFAREA 7.542800 ;
    PORT
      LAYER met4 ;
        RECT 8.000 5.000 9.200 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 34.580 167.925 39.810 173.790 ;
        RECT 47.045 171.940 119.455 188.360 ;
        RECT 34.580 165.935 45.535 167.925 ;
        RECT 34.580 165.925 39.810 165.935 ;
        RECT 47.045 165.820 81.145 171.940 ;
      LAYER pwell ;
        RECT 95.800 169.835 97.300 171.095 ;
        RECT 38.060 165.590 39.750 165.620 ;
        RECT 34.630 165.330 40.310 165.590 ;
        RECT 34.630 165.160 40.490 165.330 ;
        RECT 34.630 159.790 35.060 165.160 ;
        RECT 34.140 159.360 35.060 159.790 ;
        RECT 34.140 158.125 34.570 159.360 ;
        RECT 35.580 158.420 36.340 165.010 ;
        RECT 39.880 164.900 40.490 165.160 ;
        RECT 34.140 157.695 37.100 158.125 ;
        RECT 36.670 154.970 37.100 157.695 ;
        RECT 36.525 154.540 37.100 154.970 ;
        RECT 36.525 153.545 36.955 154.540 ;
        RECT 37.250 153.840 39.910 164.740 ;
        RECT 40.060 154.970 40.490 164.900 ;
        RECT 40.640 163.685 41.940 165.585 ;
        RECT 42.110 163.685 43.050 165.585 ;
        RECT 43.080 163.685 44.450 165.585 ;
        RECT 44.545 163.685 45.485 165.585 ;
        RECT 47.040 164.890 82.010 165.320 ;
        RECT 47.040 158.060 72.020 164.890 ;
        RECT 72.030 161.610 75.320 164.370 ;
        RECT 75.340 161.610 81.410 164.370 ;
        RECT 72.030 158.200 75.320 161.600 ;
        RECT 75.340 158.200 81.410 161.600 ;
        RECT 81.580 158.060 82.010 164.890 ;
        RECT 47.040 157.630 82.010 158.060 ;
        RECT 47.040 156.840 56.510 157.630 ;
        RECT 47.040 155.530 47.470 156.840 ;
        RECT 56.080 155.530 56.510 156.840 ;
        RECT 40.060 154.540 40.635 154.970 ;
        RECT 40.205 153.545 40.635 154.540 ;
        RECT 36.525 153.115 40.635 153.545 ;
        RECT 47.040 147.050 56.510 155.530 ;
        RECT 57.480 155.395 58.740 156.895 ;
        RECT 63.210 156.600 73.230 157.630 ;
        RECT 63.210 155.550 63.640 156.600 ;
        RECT 72.800 155.550 73.230 156.600 ;
        RECT 63.210 155.120 73.230 155.550 ;
        RECT 35.780 142.245 55.360 143.010 ;
        RECT 35.780 137.075 36.545 142.245 ;
        RECT 41.715 137.075 42.985 142.245 ;
        RECT 48.155 137.075 49.425 142.245 ;
        RECT 54.595 137.075 55.360 142.245 ;
        RECT 35.780 135.805 55.360 137.075 ;
        RECT 35.780 130.635 36.545 135.805 ;
        RECT 41.715 130.635 42.985 135.805 ;
        RECT 48.155 130.635 49.425 135.805 ;
        RECT 54.595 130.635 55.360 135.805 ;
        RECT 35.780 129.365 55.360 130.635 ;
        RECT 35.780 124.195 36.545 129.365 ;
        RECT 41.715 124.195 42.985 129.365 ;
        RECT 48.155 124.195 49.425 129.365 ;
        RECT 54.595 124.195 55.360 129.365 ;
        RECT 35.780 123.430 55.360 124.195 ;
      LAYER nwell ;
        RECT 44.640 76.045 49.870 81.910 ;
        RECT 57.105 80.060 129.515 96.480 ;
        RECT 44.640 74.055 55.595 76.045 ;
        RECT 44.640 74.045 49.870 74.055 ;
        RECT 57.105 73.940 91.205 80.060 ;
      LAYER pwell ;
        RECT 105.860 77.955 107.360 79.215 ;
        RECT 48.120 73.710 49.810 73.740 ;
        RECT 44.690 73.450 50.370 73.710 ;
        RECT 44.690 73.280 50.550 73.450 ;
        RECT 44.690 67.910 45.120 73.280 ;
        RECT 44.200 67.480 45.120 67.910 ;
        RECT 44.200 66.245 44.630 67.480 ;
        RECT 45.640 66.540 46.400 73.130 ;
        RECT 49.940 73.020 50.550 73.280 ;
        RECT 44.200 65.815 47.160 66.245 ;
        RECT 46.730 63.090 47.160 65.815 ;
        RECT 46.585 62.660 47.160 63.090 ;
        RECT 46.585 61.665 47.015 62.660 ;
        RECT 47.310 61.960 49.970 72.860 ;
        RECT 50.120 63.090 50.550 73.020 ;
        RECT 50.700 71.805 52.000 73.705 ;
        RECT 52.170 71.805 53.110 73.705 ;
        RECT 53.140 71.805 54.510 73.705 ;
        RECT 54.605 71.805 55.545 73.705 ;
        RECT 57.100 73.010 92.070 73.440 ;
        RECT 50.120 62.660 50.695 63.090 ;
        RECT 50.265 61.665 50.695 62.660 ;
        RECT 46.585 61.235 50.695 61.665 ;
        RECT 57.100 55.600 57.530 73.010 ;
        RECT 58.035 64.960 65.665 72.860 ;
        RECT 66.140 66.180 67.010 73.010 ;
        RECT 67.140 69.730 75.990 72.490 ;
        RECT 76.010 69.730 82.080 72.490 ;
        RECT 82.090 69.730 85.380 72.490 ;
        RECT 85.400 69.730 91.470 72.490 ;
        RECT 67.140 66.320 75.990 69.720 ;
        RECT 76.010 66.320 82.080 69.720 ;
        RECT 82.090 66.320 85.380 69.720 ;
        RECT 85.400 66.320 91.470 69.720 ;
        RECT 91.640 66.180 92.070 73.010 ;
        RECT 66.140 65.750 92.070 66.180 ;
        RECT 58.035 55.750 65.665 63.650 ;
        RECT 66.140 55.600 66.570 65.750 ;
        RECT 67.540 63.515 68.800 65.015 ;
        RECT 73.270 64.720 83.290 65.150 ;
        RECT 73.270 63.670 73.700 64.720 ;
        RECT 82.860 63.670 83.290 64.720 ;
        RECT 73.270 63.240 83.290 63.670 ;
        RECT 57.100 55.170 66.570 55.600 ;
        RECT 45.840 50.365 65.420 51.130 ;
        RECT 45.840 45.195 46.605 50.365 ;
        RECT 51.775 45.195 53.045 50.365 ;
        RECT 58.215 45.195 59.485 50.365 ;
        RECT 64.655 45.195 65.420 50.365 ;
        RECT 45.840 43.925 65.420 45.195 ;
        RECT 45.840 38.755 46.605 43.925 ;
        RECT 51.775 38.755 53.045 43.925 ;
        RECT 58.215 38.755 59.485 43.925 ;
        RECT 64.655 38.755 65.420 43.925 ;
        RECT 45.840 37.485 65.420 38.755 ;
        RECT 45.840 32.315 46.605 37.485 ;
        RECT 51.775 32.315 53.045 37.485 ;
        RECT 58.215 32.315 59.485 37.485 ;
        RECT 64.655 32.315 65.420 37.485 ;
        RECT 45.840 31.550 65.420 32.315 ;
      LAYER li1 ;
        RECT 47.225 188.010 119.275 188.180 ;
        RECT 47.225 187.550 47.395 188.010 ;
        RECT 75.845 187.550 76.545 188.010 ;
        RECT 47.225 187.460 76.545 187.550 ;
        RECT 90.915 187.460 91.615 188.010 ;
        RECT 119.105 187.460 119.275 188.010 ;
        RECT 47.225 187.280 119.275 187.460 ;
        RECT 28.020 178.760 28.370 180.920 ;
        RECT 28.580 178.760 28.930 180.920 ;
        RECT 29.140 178.760 29.490 180.920 ;
        RECT 29.700 178.760 30.050 180.920 ;
        RECT 30.260 178.760 30.610 180.920 ;
        RECT 30.820 178.760 31.170 180.920 ;
        RECT 31.380 178.760 31.730 180.920 ;
        RECT 31.940 178.760 32.290 180.920 ;
        RECT 32.500 178.760 32.850 180.920 ;
        RECT 33.060 178.760 33.410 180.920 ;
        RECT 34.760 173.440 39.630 173.610 ;
        RECT 34.760 167.960 34.930 173.440 ;
        RECT 39.460 172.985 39.630 173.440 ;
        RECT 38.895 172.980 39.630 172.985 ;
        RECT 37.260 172.535 39.630 172.980 ;
        RECT 37.260 172.530 39.010 172.535 ;
        RECT 37.260 172.045 37.810 172.530 ;
        RECT 38.460 172.045 39.010 172.530 ;
        RECT 34.760 167.680 36.710 167.960 ;
        RECT 34.760 166.275 34.930 167.680 ;
        RECT 35.270 166.900 35.500 167.230 ;
        RECT 35.710 167.195 36.710 167.680 ;
        RECT 38.020 166.935 38.250 171.990 ;
        RECT 39.460 167.685 39.630 172.535 ;
        RECT 47.225 172.290 47.395 187.280 ;
        RECT 47.885 173.070 48.055 186.930 ;
        RECT 51.165 173.070 51.335 186.930 ;
        RECT 51.695 174.985 51.865 186.930 ;
        RECT 54.975 182.900 55.145 186.930 ;
        RECT 58.250 186.910 58.430 187.280 ;
        RECT 54.975 181.850 55.150 182.900 ;
        RECT 51.695 174.815 51.875 174.985 ;
        RECT 51.695 173.070 51.865 174.815 ;
        RECT 54.975 173.070 55.145 181.850 ;
        RECT 58.255 173.070 58.425 186.910 ;
        RECT 61.535 173.070 61.705 186.930 ;
        RECT 64.810 186.900 64.990 187.280 ;
        RECT 75.845 187.190 119.275 187.280 ;
        RECT 64.815 173.070 64.985 186.900 ;
        RECT 68.095 182.900 68.265 186.930 ;
        RECT 68.090 181.850 68.265 182.900 ;
        RECT 68.095 173.070 68.265 181.850 ;
        RECT 71.375 174.985 71.545 186.930 ;
        RECT 71.365 174.815 71.545 174.985 ;
        RECT 71.375 173.070 71.545 174.815 ;
        RECT 71.905 173.070 72.075 186.930 ;
        RECT 75.185 173.070 75.355 186.930 ;
        RECT 48.110 172.630 51.110 172.860 ;
        RECT 51.920 172.630 54.920 172.860 ;
        RECT 55.200 172.630 58.200 172.860 ;
        RECT 58.480 172.630 61.480 172.860 ;
        RECT 61.760 172.630 64.760 172.860 ;
        RECT 65.040 172.630 68.040 172.860 ;
        RECT 68.320 172.630 71.320 172.860 ;
        RECT 72.130 172.630 75.130 172.860 ;
        RECT 75.845 172.290 76.545 187.190 ;
        RECT 77.085 173.070 77.255 186.840 ;
        RECT 80.365 173.070 80.535 186.840 ;
        RECT 83.640 186.820 83.820 187.190 ;
        RECT 83.645 173.070 83.815 186.820 ;
        RECT 86.925 173.070 87.095 186.840 ;
        RECT 90.205 173.070 90.375 186.840 ;
        RECT 77.310 172.630 80.310 172.860 ;
        RECT 80.590 172.630 83.590 172.860 ;
        RECT 83.870 172.630 86.870 172.860 ;
        RECT 87.150 172.630 90.150 172.860 ;
        RECT 90.915 172.290 91.615 187.190 ;
        RECT 92.155 173.070 92.325 186.840 ;
        RECT 95.435 173.070 95.605 186.840 ;
        RECT 98.715 173.070 98.885 187.190 ;
        RECT 101.995 173.070 102.165 186.840 ;
        RECT 105.275 173.070 105.445 186.840 ;
        RECT 108.550 186.790 108.730 187.190 ;
        RECT 108.555 173.070 108.725 186.790 ;
        RECT 111.835 172.860 112.005 186.840 ;
        RECT 115.110 186.770 115.290 187.190 ;
        RECT 115.115 173.070 115.285 186.770 ;
        RECT 118.395 173.070 118.565 186.840 ;
        RECT 92.380 172.630 95.380 172.860 ;
        RECT 95.660 172.630 98.660 172.860 ;
        RECT 98.940 172.630 101.940 172.860 ;
        RECT 102.220 172.630 105.220 172.860 ;
        RECT 105.500 172.630 108.500 172.860 ;
        RECT 108.780 172.630 115.060 172.860 ;
        RECT 115.340 172.630 118.340 172.860 ;
        RECT 119.105 172.290 119.275 187.190 ;
        RECT 47.225 172.200 119.275 172.290 ;
        RECT 46.330 172.120 119.275 172.200 ;
        RECT 46.330 171.760 47.520 172.120 ;
        RECT 58.460 171.760 58.750 172.120 ;
        RECT 46.330 171.610 58.905 171.760 ;
        RECT 59.270 171.750 59.560 172.120 ;
        RECT 64.250 171.750 64.600 172.120 ;
        RECT 64.960 171.755 65.310 172.120 ;
        RECT 80.500 171.760 80.960 172.120 ;
        RECT 76.015 171.755 80.965 171.760 ;
        RECT 47.225 171.590 58.905 171.610 ;
        RECT 47.225 170.490 47.395 171.590 ;
        RECT 58.735 170.940 58.905 171.590 ;
        RECT 56.870 170.935 58.905 170.940 ;
        RECT 48.875 170.705 51.605 170.935 ;
        RECT 48.285 170.490 48.555 170.495 ;
        RECT 47.225 169.860 48.555 170.490 ;
        RECT 40.170 167.920 42.190 168.220 ;
        RECT 42.915 167.955 43.295 168.315 ;
        RECT 39.410 167.515 39.680 167.685 ;
        RECT 35.710 166.765 38.250 166.935 ;
        RECT 38.460 166.765 39.010 166.935 ;
        RECT 39.460 166.275 39.630 167.515 ;
        RECT 40.170 166.700 40.470 167.920 ;
        RECT 40.780 167.465 41.870 167.735 ;
        RECT 42.250 167.465 42.910 167.735 ;
        RECT 43.290 167.465 44.310 167.735 ;
        RECT 44.685 167.465 45.345 167.735 ;
        RECT 34.760 166.105 39.630 166.275 ;
        RECT 37.570 165.880 37.810 165.890 ;
        RECT 40.370 165.880 40.610 165.970 ;
        RECT 37.570 165.660 40.610 165.880 ;
        RECT 40.810 165.915 40.980 167.115 ;
        RECT 41.240 166.115 41.410 167.465 ;
        RECT 41.670 165.930 41.840 167.115 ;
        RECT 42.280 166.115 42.450 167.465 ;
        RECT 41.670 165.915 42.530 165.930 ;
        RECT 40.810 165.745 42.530 165.915 ;
        RECT 37.570 165.650 37.810 165.660 ;
        RECT 40.370 165.580 40.610 165.660 ;
        RECT 41.670 165.630 42.530 165.745 ;
        RECT 38.190 165.460 39.620 165.490 ;
        RECT 34.760 165.320 40.180 165.460 ;
        RECT 41.670 165.455 41.840 165.630 ;
        RECT 34.760 165.290 38.360 165.320 ;
        RECT 39.450 165.290 40.180 165.320 ;
        RECT 28.020 159.260 28.370 161.420 ;
        RECT 28.580 159.260 28.930 161.420 ;
        RECT 29.140 159.260 29.490 161.420 ;
        RECT 29.700 159.260 30.050 161.420 ;
        RECT 30.260 159.260 30.610 161.420 ;
        RECT 30.820 159.260 31.170 161.420 ;
        RECT 31.380 159.260 31.730 161.420 ;
        RECT 31.940 159.260 32.290 161.420 ;
        RECT 32.500 159.260 32.850 161.420 ;
        RECT 33.060 159.260 33.410 161.420 ;
        RECT 34.760 159.660 34.930 165.290 ;
        RECT 40.010 165.200 40.180 165.290 ;
        RECT 35.710 164.670 36.210 164.840 ;
        RECT 36.830 164.670 37.230 165.120 ;
        RECT 40.010 165.030 40.360 165.200 ;
        RECT 37.850 164.850 39.740 165.020 ;
        RECT 34.270 159.490 34.930 159.660 ;
        RECT 35.270 159.615 35.500 164.615 ;
        RECT 34.270 157.995 34.440 159.490 ;
        RECT 35.710 157.995 36.210 159.560 ;
        RECT 34.270 157.825 36.970 157.995 ;
        RECT 36.800 154.840 36.970 157.825 ;
        RECT 36.655 154.670 36.970 154.840 ;
        RECT 36.655 154.250 36.825 154.670 ;
        RECT 37.420 154.250 37.590 164.610 ;
        RECT 37.850 154.610 38.020 164.850 ;
        RECT 38.280 154.250 38.450 164.610 ;
        RECT 38.710 154.610 38.880 164.850 ;
        RECT 39.140 154.250 39.310 164.610 ;
        RECT 39.570 154.610 39.740 164.850 ;
        RECT 40.190 164.110 40.360 165.030 ;
        RECT 40.810 164.110 40.980 165.455 ;
        RECT 41.600 165.285 41.840 165.455 ;
        RECT 41.600 164.455 41.770 165.285 ;
        RECT 42.280 164.110 42.450 165.455 ;
        RECT 42.710 164.800 42.880 167.115 ;
        RECT 43.320 166.115 43.490 167.465 ;
        RECT 44.720 167.180 44.890 167.465 ;
        RECT 44.110 165.930 44.280 167.115 ;
        RECT 44.700 167.010 44.890 167.180 ;
        RECT 44.715 166.115 44.885 167.010 ;
        RECT 44.110 165.870 44.940 165.930 ;
        RECT 43.680 165.630 44.940 165.870 ;
        RECT 45.145 165.920 45.315 167.115 ;
        RECT 47.225 166.170 47.395 169.860 ;
        RECT 48.285 167.495 48.555 169.860 ;
        RECT 48.875 167.285 49.045 170.705 ;
        RECT 50.155 167.285 50.325 170.705 ;
        RECT 51.435 167.495 51.605 170.705 ;
        RECT 54.525 170.705 58.905 170.935 ;
        RECT 52.715 167.285 52.885 170.495 ;
        RECT 53.245 167.495 53.415 170.495 ;
        RECT 54.525 167.495 54.695 170.705 ;
        RECT 55.805 167.495 55.975 170.705 ;
        RECT 56.870 170.700 58.905 170.705 ;
        RECT 57.085 167.285 57.255 170.700 ;
        RECT 57.575 167.495 57.845 170.495 ;
        RECT 48.875 167.055 51.380 167.285 ;
        RECT 51.660 167.055 52.885 167.285 ;
        RECT 53.470 167.055 54.470 167.285 ;
        RECT 54.750 167.055 55.750 167.285 ;
        RECT 56.030 167.055 57.255 167.285 ;
        RECT 58.735 166.170 58.905 170.700 ;
        RECT 47.225 166.000 58.905 166.170 ;
        RECT 59.265 171.670 64.600 171.750 ;
        RECT 59.265 171.580 64.595 171.670 ;
        RECT 59.265 171.240 59.435 171.580 ;
        RECT 64.425 171.240 64.595 171.580 ;
        RECT 64.955 171.590 80.965 171.755 ;
        RECT 64.955 171.585 76.185 171.590 ;
        RECT 64.955 171.240 65.125 171.585 ;
        RECT 59.265 171.150 65.130 171.240 ;
        RECT 80.795 171.150 80.965 171.590 ;
        RECT 59.265 170.970 80.965 171.150 ;
        RECT 59.265 166.170 59.435 170.970 ;
        RECT 59.815 167.070 59.985 170.970 ;
        RECT 61.095 167.070 61.265 170.620 ;
        RECT 62.375 167.070 62.545 170.970 ;
        RECT 64.370 170.880 80.965 170.970 ;
        RECT 63.655 167.070 63.825 170.620 ;
        RECT 60.040 166.630 61.040 166.860 ;
        RECT 61.320 166.630 62.320 166.860 ;
        RECT 62.600 166.630 63.600 166.860 ;
        RECT 64.425 166.170 64.595 170.880 ;
        RECT 59.265 166.000 64.595 166.170 ;
        RECT 64.955 166.170 65.125 170.880 ;
        RECT 65.485 166.945 65.655 170.880 ;
        RECT 68.765 166.945 68.935 170.880 ;
        RECT 69.375 167.155 69.545 170.530 ;
        RECT 72.655 167.155 72.825 170.880 ;
        RECT 75.935 166.945 76.105 170.530 ;
        RECT 65.485 166.715 68.935 166.945 ;
        RECT 69.600 166.715 72.600 166.945 ;
        RECT 72.880 166.715 76.105 166.945 ;
        RECT 76.545 166.945 76.715 170.880 ;
        RECT 79.825 166.945 79.995 170.880 ;
        RECT 76.545 166.715 79.995 166.945 ;
        RECT 80.795 166.170 80.965 170.880 ;
        RECT 82.450 169.300 83.860 171.460 ;
        RECT 84.070 169.300 85.480 171.460 ;
        RECT 85.690 169.300 87.100 171.460 ;
        RECT 87.310 169.300 88.720 171.460 ;
        RECT 88.930 169.300 90.340 171.460 ;
        RECT 90.550 169.300 91.960 171.460 ;
        RECT 92.170 169.300 93.580 171.460 ;
        RECT 93.790 169.300 95.200 171.460 ;
        RECT 96.745 171.290 96.915 171.620 ;
        RECT 95.940 169.965 96.700 170.965 ;
        RECT 96.960 169.965 97.130 170.965 ;
        RECT 96.650 169.150 97.000 169.510 ;
        RECT 64.955 166.000 80.965 166.170 ;
        RECT 42.650 164.470 42.950 164.800 ;
        RECT 42.710 164.455 42.880 164.470 ;
        RECT 43.250 164.110 43.420 165.455 ;
        RECT 43.680 164.455 43.850 165.630 ;
        RECT 45.145 165.600 45.730 165.920 ;
        RECT 44.110 164.110 44.280 165.455 ;
        RECT 44.715 164.110 44.885 165.455 ;
        RECT 45.145 164.455 45.315 165.600 ;
        RECT 47.170 165.020 81.880 165.190 ;
        RECT 47.170 164.600 47.340 165.020 ;
        RECT 47.170 164.330 55.465 164.600 ;
        RECT 47.170 164.110 47.340 164.330 ;
        RECT 40.190 163.810 47.340 164.110 ;
        RECT 40.190 154.840 40.360 163.810 ;
        RECT 44.350 163.280 44.690 163.630 ;
        RECT 40.190 154.670 40.505 154.840 ;
        RECT 40.335 154.250 40.505 154.670 ;
        RECT 36.655 153.980 40.505 154.250 ;
        RECT 36.655 153.415 36.825 153.980 ;
        RECT 40.335 153.415 40.505 153.980 ;
        RECT 36.655 153.245 40.505 153.415 ;
        RECT 47.170 148.040 47.340 163.810 ;
        RECT 48.145 156.970 48.315 163.970 ;
        RECT 49.925 156.970 50.095 163.970 ;
        RECT 51.705 156.970 51.875 163.970 ;
        RECT 53.485 156.970 53.655 163.970 ;
        RECT 55.265 162.950 55.435 163.970 ;
        RECT 55.265 162.650 55.690 162.950 ;
        RECT 55.265 156.970 55.435 162.650 ;
        RECT 56.210 157.930 56.380 165.020 ;
        RECT 56.650 164.680 56.820 165.020 ;
        RECT 81.710 164.680 81.880 165.020 ;
        RECT 56.630 164.450 59.975 164.680 ;
        RECT 60.255 164.450 62.755 164.680 ;
        RECT 63.035 164.450 65.535 164.680 ;
        RECT 66.120 164.450 68.845 164.680 ;
        RECT 69.125 164.450 71.955 164.680 ;
        RECT 72.425 164.450 74.925 164.680 ;
        RECT 75.735 164.450 78.235 164.680 ;
        RECT 78.515 164.450 81.880 164.680 ;
        RECT 82.450 164.610 83.860 166.770 ;
        RECT 84.070 164.610 85.480 166.770 ;
        RECT 85.690 164.610 87.100 166.770 ;
        RECT 87.310 164.610 88.720 166.770 ;
        RECT 88.930 164.610 90.340 166.770 ;
        RECT 90.550 164.610 91.960 166.770 ;
        RECT 92.170 164.610 93.580 166.770 ;
        RECT 93.790 164.610 95.200 166.770 ;
        RECT 96.090 166.480 97.500 168.640 ;
        RECT 97.710 166.480 99.120 168.640 ;
        RECT 99.330 166.480 100.740 168.640 ;
        RECT 100.950 166.480 102.360 168.640 ;
        RECT 102.570 166.480 103.980 168.640 ;
        RECT 104.190 166.480 105.600 168.640 ;
        RECT 105.810 166.480 107.220 168.640 ;
        RECT 107.430 166.480 108.840 168.640 ;
        RECT 109.180 166.880 111.340 168.290 ;
        RECT 116.780 166.880 118.940 168.290 ;
        RECT 109.180 165.230 111.340 166.640 ;
        RECT 116.780 165.230 118.940 166.640 ;
        RECT 56.650 158.610 56.820 164.450 ;
        RECT 57.250 158.610 57.420 164.450 ;
        RECT 60.030 158.610 60.200 164.240 ;
        RECT 62.810 158.970 62.980 164.240 ;
        RECT 65.590 158.610 65.760 164.240 ;
        RECT 66.120 158.970 66.290 164.450 ;
        RECT 68.900 158.610 69.070 164.240 ;
        RECT 71.680 158.970 71.850 164.450 ;
        RECT 72.200 158.610 72.370 164.240 ;
        RECT 74.980 158.970 75.150 164.240 ;
        RECT 75.510 158.970 75.680 164.240 ;
        RECT 78.290 158.610 78.460 164.240 ;
        RECT 81.070 158.610 81.240 164.450 ;
        RECT 81.710 158.610 81.880 164.450 ;
        RECT 82.450 162.240 83.860 164.400 ;
        RECT 84.070 162.240 85.480 164.400 ;
        RECT 85.690 162.240 87.100 164.400 ;
        RECT 87.310 162.240 88.720 164.400 ;
        RECT 88.930 162.240 90.340 164.400 ;
        RECT 90.550 162.240 91.960 164.400 ;
        RECT 92.170 162.240 93.580 164.400 ;
        RECT 93.790 162.240 95.200 164.400 ;
        RECT 96.090 162.120 97.500 164.280 ;
        RECT 97.710 162.120 99.120 164.280 ;
        RECT 99.330 162.120 100.740 164.280 ;
        RECT 100.950 162.120 102.360 164.280 ;
        RECT 102.570 162.120 103.980 164.280 ;
        RECT 104.190 162.120 105.600 164.280 ;
        RECT 105.810 162.120 107.220 164.280 ;
        RECT 107.430 162.120 108.840 164.280 ;
        RECT 109.180 163.580 111.340 164.990 ;
        RECT 116.780 163.580 118.940 164.990 ;
        RECT 109.180 161.920 111.340 163.330 ;
        RECT 116.780 161.920 118.940 163.330 ;
        RECT 109.180 160.280 111.340 161.690 ;
        RECT 116.780 160.280 118.940 161.690 ;
        RECT 56.650 158.340 81.880 158.610 ;
        RECT 56.650 157.930 56.820 158.340 ;
        RECT 63.340 157.930 73.280 157.940 ;
        RECT 81.710 157.930 81.880 158.340 ;
        RECT 56.210 157.760 81.880 157.930 ;
        RECT 48.370 156.530 49.870 156.760 ;
        RECT 50.150 156.530 51.650 156.760 ;
        RECT 51.930 156.530 53.430 156.760 ;
        RECT 53.710 156.530 55.210 156.760 ;
        RECT 48.370 155.610 49.870 155.840 ;
        RECT 50.150 155.610 51.650 155.840 ;
        RECT 51.930 155.610 53.430 155.840 ;
        RECT 53.710 155.610 55.210 155.840 ;
        RECT 48.145 148.400 48.315 155.400 ;
        RECT 49.925 150.770 50.095 155.400 ;
        RECT 49.920 149.000 50.100 150.770 ;
        RECT 49.925 148.400 50.095 149.000 ;
        RECT 51.705 148.400 51.875 155.400 ;
        RECT 53.485 148.400 53.655 155.400 ;
        RECT 55.265 148.400 55.435 155.400 ;
        RECT 56.210 148.040 56.380 157.760 ;
        RECT 57.610 156.485 58.610 157.760 ;
        RECT 63.340 156.740 73.280 157.760 ;
        RECT 82.450 157.550 83.860 159.710 ;
        RECT 84.070 157.550 85.480 159.710 ;
        RECT 85.690 157.550 87.100 159.710 ;
        RECT 87.310 157.550 88.720 159.710 ;
        RECT 88.930 157.550 90.340 159.710 ;
        RECT 90.550 157.550 91.960 159.710 ;
        RECT 92.170 157.550 93.580 159.710 ;
        RECT 93.790 157.550 95.200 159.710 ;
        RECT 109.180 158.630 111.340 160.040 ;
        RECT 116.780 158.630 118.940 160.040 ;
        RECT 109.180 156.980 111.340 158.390 ;
        RECT 116.780 156.980 118.940 158.390 ;
        RECT 63.340 156.730 73.100 156.740 ;
        RECT 56.880 155.690 57.230 156.030 ;
        RECT 57.610 155.995 59.500 156.165 ;
        RECT 57.610 155.565 58.610 155.735 ;
        RECT 63.340 155.420 63.510 156.730 ;
        RECT 63.990 155.900 66.150 156.250 ;
        RECT 70.290 155.900 72.450 156.250 ;
        RECT 72.930 155.420 73.100 156.730 ;
        RECT 63.340 155.250 73.100 155.420 ;
        RECT 109.180 155.330 111.340 156.740 ;
        RECT 116.780 155.330 118.940 156.740 ;
        RECT 57.430 152.440 58.840 154.600 ;
        RECT 59.080 152.440 60.490 154.600 ;
        RECT 64.980 152.440 66.390 154.600 ;
        RECT 66.630 152.440 68.040 154.600 ;
        RECT 47.170 147.770 56.380 148.040 ;
        RECT 47.170 147.350 47.340 147.770 ;
        RECT 56.210 147.350 56.380 147.770 ;
        RECT 47.170 147.180 56.380 147.350 ;
        RECT 47.170 142.880 48.200 147.180 ;
        RECT 61.180 144.370 64.290 146.530 ;
        RECT 35.910 142.385 55.230 142.880 ;
        RECT 35.910 136.935 36.405 142.385 ;
        RECT 36.725 141.705 41.535 142.065 ;
        RECT 36.725 137.615 37.085 141.705 ;
        RECT 37.395 137.925 40.865 141.395 ;
        RECT 41.175 137.615 41.535 141.705 ;
        RECT 36.725 137.255 41.535 137.615 ;
        RECT 41.180 136.935 41.530 137.255 ;
        RECT 41.855 136.935 42.845 142.385 ;
        RECT 43.165 141.705 47.975 142.065 ;
        RECT 43.165 137.615 43.525 141.705 ;
        RECT 43.835 137.925 47.305 141.395 ;
        RECT 47.615 137.615 47.975 141.705 ;
        RECT 43.165 137.255 47.975 137.615 ;
        RECT 43.170 136.935 43.520 137.255 ;
        RECT 47.620 136.935 47.970 137.255 ;
        RECT 48.295 136.935 49.285 142.385 ;
        RECT 49.605 141.705 54.415 142.065 ;
        RECT 49.605 137.615 49.965 141.705 ;
        RECT 50.275 137.925 53.745 141.395 ;
        RECT 54.055 137.940 54.415 141.705 ;
        RECT 54.055 137.615 54.420 137.940 ;
        RECT 49.605 137.255 54.420 137.615 ;
        RECT 49.610 136.935 49.960 137.255 ;
        RECT 54.070 136.935 54.420 137.255 ;
        RECT 54.735 136.935 55.230 142.385 ;
        RECT 61.180 137.170 62.590 142.240 ;
        RECT 62.880 140.080 64.290 142.240 ;
        RECT 62.880 137.170 64.290 139.330 ;
        RECT 35.910 135.945 55.230 136.935 ;
        RECT 35.910 130.495 36.405 135.945 ;
        RECT 41.180 135.625 41.530 135.945 ;
        RECT 36.725 135.265 41.535 135.625 ;
        RECT 36.725 131.175 37.085 135.265 ;
        RECT 37.395 131.485 40.865 134.955 ;
        RECT 41.175 131.175 41.535 135.265 ;
        RECT 36.725 130.815 41.535 131.175 ;
        RECT 41.180 130.495 41.530 130.815 ;
        RECT 41.855 130.495 42.845 135.945 ;
        RECT 43.170 135.625 43.520 135.945 ;
        RECT 47.620 135.625 47.970 135.945 ;
        RECT 43.165 135.265 47.975 135.625 ;
        RECT 43.165 131.175 43.525 135.265 ;
        RECT 43.835 131.485 47.305 134.955 ;
        RECT 47.615 131.175 47.975 135.265 ;
        RECT 43.165 130.815 47.975 131.175 ;
        RECT 43.170 130.495 43.520 130.815 ;
        RECT 47.620 130.495 47.970 130.815 ;
        RECT 48.295 130.495 49.285 135.945 ;
        RECT 49.610 135.625 49.960 135.945 ;
        RECT 54.070 135.625 54.420 135.945 ;
        RECT 49.605 135.265 54.420 135.625 ;
        RECT 49.605 131.175 49.965 135.265 ;
        RECT 50.275 131.485 53.745 134.955 ;
        RECT 54.055 131.175 54.420 135.265 ;
        RECT 49.605 130.815 54.420 131.175 ;
        RECT 49.610 130.495 49.960 130.815 ;
        RECT 54.070 130.495 54.420 130.815 ;
        RECT 54.735 130.495 55.230 135.945 ;
        RECT 61.180 132.880 64.290 135.040 ;
        RECT 35.910 129.505 55.230 130.495 ;
        RECT 35.910 124.055 36.405 129.505 ;
        RECT 41.180 129.185 41.530 129.505 ;
        RECT 36.725 128.825 41.535 129.185 ;
        RECT 36.725 124.735 37.085 128.825 ;
        RECT 37.395 125.045 40.865 128.515 ;
        RECT 41.175 124.735 41.535 128.825 ;
        RECT 36.725 124.375 41.535 124.735 ;
        RECT 41.855 124.055 42.845 129.505 ;
        RECT 43.170 129.185 43.520 129.505 ;
        RECT 47.620 129.185 47.970 129.505 ;
        RECT 43.165 128.825 47.975 129.185 ;
        RECT 43.165 124.735 43.525 128.825 ;
        RECT 43.835 125.045 47.305 128.515 ;
        RECT 47.615 124.735 47.975 128.825 ;
        RECT 43.165 124.375 47.975 124.735 ;
        RECT 48.295 124.055 49.285 129.505 ;
        RECT 49.610 129.185 49.960 129.505 ;
        RECT 54.070 129.185 54.420 129.505 ;
        RECT 49.605 128.830 54.420 129.185 ;
        RECT 49.605 128.825 54.415 128.830 ;
        RECT 49.605 124.735 49.965 128.825 ;
        RECT 50.275 125.045 53.745 128.515 ;
        RECT 54.055 124.735 54.415 128.825 ;
        RECT 49.605 124.375 54.415 124.735 ;
        RECT 54.735 127.900 55.230 129.505 ;
        RECT 57.430 129.330 58.840 131.490 ;
        RECT 59.080 129.330 60.490 131.490 ;
        RECT 64.980 129.330 66.390 131.490 ;
        RECT 66.630 129.330 68.040 131.490 ;
        RECT 54.735 125.740 58.840 127.900 ;
        RECT 59.080 125.740 60.490 127.900 ;
        RECT 64.980 125.740 66.390 127.900 ;
        RECT 54.735 124.060 55.230 125.740 ;
        RECT 66.630 124.060 68.040 127.900 ;
        RECT 54.620 124.055 68.040 124.060 ;
        RECT 35.910 123.560 68.040 124.055 ;
        RECT 57.430 102.630 58.840 104.790 ;
        RECT 59.080 102.630 60.490 104.790 ;
        RECT 64.980 102.630 66.390 104.790 ;
        RECT 66.630 102.630 68.040 104.790 ;
        RECT 57.285 96.130 129.335 96.300 ;
        RECT 57.285 95.670 57.455 96.130 ;
        RECT 85.905 95.670 86.605 96.130 ;
        RECT 57.285 95.580 86.605 95.670 ;
        RECT 100.975 95.580 101.675 96.130 ;
        RECT 129.165 95.580 129.335 96.130 ;
        RECT 57.285 95.400 129.335 95.580 ;
        RECT 38.080 86.880 38.430 89.040 ;
        RECT 38.640 86.880 38.990 89.040 ;
        RECT 39.200 86.880 39.550 89.040 ;
        RECT 39.760 86.880 40.110 89.040 ;
        RECT 40.320 86.880 40.670 89.040 ;
        RECT 40.880 86.880 41.230 89.040 ;
        RECT 41.440 86.880 41.790 89.040 ;
        RECT 42.000 86.880 42.350 89.040 ;
        RECT 42.560 86.880 42.910 89.040 ;
        RECT 43.120 86.880 43.470 89.040 ;
        RECT 44.820 81.560 49.690 81.730 ;
        RECT 44.820 76.080 44.990 81.560 ;
        RECT 49.520 81.105 49.690 81.560 ;
        RECT 48.955 81.100 49.690 81.105 ;
        RECT 47.320 80.655 49.690 81.100 ;
        RECT 47.320 80.650 49.070 80.655 ;
        RECT 47.320 80.165 47.870 80.650 ;
        RECT 48.520 80.165 49.070 80.650 ;
        RECT 44.820 75.800 46.770 76.080 ;
        RECT 44.820 74.395 44.990 75.800 ;
        RECT 45.330 75.020 45.560 75.350 ;
        RECT 45.770 75.315 46.770 75.800 ;
        RECT 48.080 75.055 48.310 80.110 ;
        RECT 49.520 75.805 49.690 80.655 ;
        RECT 57.285 80.410 57.455 95.400 ;
        RECT 57.945 81.190 58.115 95.050 ;
        RECT 61.225 81.190 61.395 95.050 ;
        RECT 61.755 83.105 61.925 95.050 ;
        RECT 65.035 91.020 65.205 95.050 ;
        RECT 68.310 95.030 68.490 95.400 ;
        RECT 65.035 89.970 65.210 91.020 ;
        RECT 61.755 82.935 61.935 83.105 ;
        RECT 61.755 81.190 61.925 82.935 ;
        RECT 65.035 81.190 65.205 89.970 ;
        RECT 68.315 81.190 68.485 95.030 ;
        RECT 71.595 81.190 71.765 95.050 ;
        RECT 74.870 95.020 75.050 95.400 ;
        RECT 85.905 95.310 129.335 95.400 ;
        RECT 74.875 81.190 75.045 95.020 ;
        RECT 78.155 91.020 78.325 95.050 ;
        RECT 78.150 89.970 78.325 91.020 ;
        RECT 78.155 81.190 78.325 89.970 ;
        RECT 81.435 83.105 81.605 95.050 ;
        RECT 81.425 82.935 81.605 83.105 ;
        RECT 81.435 81.190 81.605 82.935 ;
        RECT 81.965 81.190 82.135 95.050 ;
        RECT 85.245 81.190 85.415 95.050 ;
        RECT 58.170 80.750 61.170 80.980 ;
        RECT 61.980 80.750 64.980 80.980 ;
        RECT 65.260 80.750 68.260 80.980 ;
        RECT 68.540 80.750 71.540 80.980 ;
        RECT 71.820 80.750 74.820 80.980 ;
        RECT 75.100 80.750 78.100 80.980 ;
        RECT 78.380 80.750 81.380 80.980 ;
        RECT 82.190 80.750 85.190 80.980 ;
        RECT 85.905 80.410 86.605 95.310 ;
        RECT 87.145 81.190 87.315 94.960 ;
        RECT 90.425 81.190 90.595 94.960 ;
        RECT 93.700 94.940 93.880 95.310 ;
        RECT 93.705 81.190 93.875 94.940 ;
        RECT 96.985 81.190 97.155 94.960 ;
        RECT 100.265 81.190 100.435 94.960 ;
        RECT 87.370 80.750 90.370 80.980 ;
        RECT 90.650 80.750 93.650 80.980 ;
        RECT 93.930 80.750 96.930 80.980 ;
        RECT 97.210 80.750 100.210 80.980 ;
        RECT 100.975 80.410 101.675 95.310 ;
        RECT 102.215 81.190 102.385 94.960 ;
        RECT 105.495 81.190 105.665 94.960 ;
        RECT 108.775 81.190 108.945 95.310 ;
        RECT 112.055 81.190 112.225 94.960 ;
        RECT 115.335 81.190 115.505 94.960 ;
        RECT 118.610 94.910 118.790 95.310 ;
        RECT 118.615 81.190 118.785 94.910 ;
        RECT 121.895 80.980 122.065 94.960 ;
        RECT 125.170 94.890 125.350 95.310 ;
        RECT 125.175 81.190 125.345 94.890 ;
        RECT 128.455 81.190 128.625 94.960 ;
        RECT 102.440 80.750 105.440 80.980 ;
        RECT 105.720 80.750 108.720 80.980 ;
        RECT 109.000 80.750 112.000 80.980 ;
        RECT 112.280 80.750 115.280 80.980 ;
        RECT 115.560 80.750 118.560 80.980 ;
        RECT 118.840 80.750 125.120 80.980 ;
        RECT 125.400 80.750 128.400 80.980 ;
        RECT 129.165 80.410 129.335 95.310 ;
        RECT 57.285 80.240 129.335 80.410 ;
        RECT 57.290 79.880 57.580 80.240 ;
        RECT 68.520 79.880 68.810 80.240 ;
        RECT 57.285 79.710 68.965 79.880 ;
        RECT 69.330 79.870 69.620 80.240 ;
        RECT 74.310 79.870 74.660 80.240 ;
        RECT 75.020 79.875 75.370 80.240 ;
        RECT 90.560 79.880 91.020 80.240 ;
        RECT 86.075 79.875 91.025 79.880 ;
        RECT 57.285 78.610 57.455 79.710 ;
        RECT 68.795 79.060 68.965 79.710 ;
        RECT 66.930 79.055 68.965 79.060 ;
        RECT 58.935 78.825 61.665 79.055 ;
        RECT 58.345 78.610 58.615 78.615 ;
        RECT 57.285 77.980 58.615 78.610 ;
        RECT 50.230 76.040 52.250 76.340 ;
        RECT 52.975 76.075 53.355 76.435 ;
        RECT 49.470 75.635 49.740 75.805 ;
        RECT 45.770 74.885 48.310 75.055 ;
        RECT 48.520 74.885 49.070 75.055 ;
        RECT 49.520 74.395 49.690 75.635 ;
        RECT 50.230 74.820 50.530 76.040 ;
        RECT 50.840 75.585 51.930 75.855 ;
        RECT 52.310 75.585 52.970 75.855 ;
        RECT 53.350 75.585 54.370 75.855 ;
        RECT 54.745 75.585 55.405 75.855 ;
        RECT 44.820 74.225 49.690 74.395 ;
        RECT 47.630 74.000 47.870 74.010 ;
        RECT 50.430 74.000 50.670 74.090 ;
        RECT 47.630 73.780 50.670 74.000 ;
        RECT 50.870 74.035 51.040 75.235 ;
        RECT 51.300 74.235 51.470 75.585 ;
        RECT 51.730 74.050 51.900 75.235 ;
        RECT 52.340 74.235 52.510 75.585 ;
        RECT 51.730 74.035 52.590 74.050 ;
        RECT 50.870 73.865 52.590 74.035 ;
        RECT 47.630 73.770 47.870 73.780 ;
        RECT 50.430 73.700 50.670 73.780 ;
        RECT 51.730 73.750 52.590 73.865 ;
        RECT 48.250 73.580 49.680 73.610 ;
        RECT 44.820 73.440 50.240 73.580 ;
        RECT 51.730 73.575 51.900 73.750 ;
        RECT 44.820 73.410 48.420 73.440 ;
        RECT 49.510 73.410 50.240 73.440 ;
        RECT 38.080 67.380 38.430 69.540 ;
        RECT 38.640 67.380 38.990 69.540 ;
        RECT 39.200 67.380 39.550 69.540 ;
        RECT 39.760 67.380 40.110 69.540 ;
        RECT 40.320 67.380 40.670 69.540 ;
        RECT 40.880 67.380 41.230 69.540 ;
        RECT 41.440 67.380 41.790 69.540 ;
        RECT 42.000 67.380 42.350 69.540 ;
        RECT 42.560 67.380 42.910 69.540 ;
        RECT 43.120 67.380 43.470 69.540 ;
        RECT 44.820 67.780 44.990 73.410 ;
        RECT 50.070 73.320 50.240 73.410 ;
        RECT 45.770 72.790 46.270 72.960 ;
        RECT 46.890 72.790 47.290 73.240 ;
        RECT 50.070 73.150 50.420 73.320 ;
        RECT 47.910 72.970 49.800 73.140 ;
        RECT 44.330 67.610 44.990 67.780 ;
        RECT 45.330 67.735 45.560 72.735 ;
        RECT 44.330 66.115 44.500 67.610 ;
        RECT 45.770 66.115 46.270 67.680 ;
        RECT 44.330 65.945 47.030 66.115 ;
        RECT 46.860 62.960 47.030 65.945 ;
        RECT 46.715 62.790 47.030 62.960 ;
        RECT 46.715 62.670 46.885 62.790 ;
        RECT 45.640 62.370 46.885 62.670 ;
        RECT 47.480 62.370 47.650 72.730 ;
        RECT 47.910 62.730 48.080 72.970 ;
        RECT 48.340 62.370 48.510 72.730 ;
        RECT 48.770 62.730 48.940 72.970 ;
        RECT 49.200 62.370 49.370 72.730 ;
        RECT 49.630 62.730 49.800 72.970 ;
        RECT 50.250 72.230 50.420 73.150 ;
        RECT 50.870 72.230 51.040 73.575 ;
        RECT 51.660 73.405 51.900 73.575 ;
        RECT 51.660 72.575 51.830 73.405 ;
        RECT 52.340 72.230 52.510 73.575 ;
        RECT 52.770 72.920 52.940 75.235 ;
        RECT 53.380 74.235 53.550 75.585 ;
        RECT 54.780 75.235 54.950 75.585 ;
        RECT 54.170 74.050 54.340 75.235 ;
        RECT 54.775 75.135 54.950 75.235 ;
        RECT 54.775 74.235 54.945 75.135 ;
        RECT 54.170 73.990 55.000 74.050 ;
        RECT 53.740 73.750 55.000 73.990 ;
        RECT 55.205 74.040 55.375 75.235 ;
        RECT 57.285 74.290 57.455 77.980 ;
        RECT 58.345 75.615 58.615 77.980 ;
        RECT 58.935 75.405 59.105 78.825 ;
        RECT 60.215 75.405 60.385 78.825 ;
        RECT 61.495 75.615 61.665 78.825 ;
        RECT 64.585 78.825 68.965 79.055 ;
        RECT 62.775 75.405 62.945 78.615 ;
        RECT 63.305 75.615 63.475 78.615 ;
        RECT 64.585 75.615 64.755 78.825 ;
        RECT 65.865 75.615 66.035 78.825 ;
        RECT 66.930 78.820 68.965 78.825 ;
        RECT 67.145 75.405 67.315 78.820 ;
        RECT 67.635 75.615 67.905 78.615 ;
        RECT 58.935 75.175 61.440 75.405 ;
        RECT 61.720 75.175 62.945 75.405 ;
        RECT 63.530 75.175 64.530 75.405 ;
        RECT 64.810 75.175 65.810 75.405 ;
        RECT 66.090 75.175 67.315 75.405 ;
        RECT 68.795 74.290 68.965 78.820 ;
        RECT 57.285 74.120 68.965 74.290 ;
        RECT 69.325 79.790 74.660 79.870 ;
        RECT 69.325 79.700 74.655 79.790 ;
        RECT 69.325 79.360 69.495 79.700 ;
        RECT 74.485 79.360 74.655 79.700 ;
        RECT 75.015 79.710 91.025 79.875 ;
        RECT 75.015 79.705 86.245 79.710 ;
        RECT 75.015 79.360 75.185 79.705 ;
        RECT 69.325 79.270 75.190 79.360 ;
        RECT 90.855 79.270 91.025 79.710 ;
        RECT 106.805 79.410 106.975 79.740 ;
        RECT 69.325 79.090 91.025 79.270 ;
        RECT 69.325 74.290 69.495 79.090 ;
        RECT 69.875 75.190 70.045 79.090 ;
        RECT 71.155 75.190 71.325 78.740 ;
        RECT 72.435 75.190 72.605 79.090 ;
        RECT 74.430 79.000 91.025 79.090 ;
        RECT 73.715 75.190 73.885 78.740 ;
        RECT 70.100 74.750 71.100 74.980 ;
        RECT 71.380 74.750 72.380 74.980 ;
        RECT 72.660 74.750 73.660 74.980 ;
        RECT 74.485 74.290 74.655 79.000 ;
        RECT 69.325 74.120 74.655 74.290 ;
        RECT 75.015 74.290 75.185 79.000 ;
        RECT 75.545 75.065 75.715 79.000 ;
        RECT 78.825 75.065 78.995 79.000 ;
        RECT 79.435 75.275 79.605 78.650 ;
        RECT 82.715 75.275 82.885 79.000 ;
        RECT 85.995 75.065 86.165 78.650 ;
        RECT 75.545 74.835 78.995 75.065 ;
        RECT 79.660 74.835 82.660 75.065 ;
        RECT 82.940 74.835 86.165 75.065 ;
        RECT 86.605 75.065 86.775 79.000 ;
        RECT 89.885 75.065 90.055 79.000 ;
        RECT 86.605 74.835 90.055 75.065 ;
        RECT 90.855 74.290 91.025 79.000 ;
        RECT 92.520 77.080 93.930 79.240 ;
        RECT 94.140 77.080 95.550 79.240 ;
        RECT 95.760 77.080 97.170 79.240 ;
        RECT 97.390 76.950 98.800 79.110 ;
        RECT 99.010 76.950 100.420 79.110 ;
        RECT 100.630 76.950 102.040 79.110 ;
        RECT 102.250 76.950 103.660 79.110 ;
        RECT 103.870 76.950 105.280 79.110 ;
        RECT 106.000 78.085 106.760 79.085 ;
        RECT 107.020 78.085 107.190 79.085 ;
        RECT 106.710 77.270 107.060 77.630 ;
        RECT 106.150 74.600 107.560 76.760 ;
        RECT 107.770 74.600 109.180 76.760 ;
        RECT 109.390 74.600 110.800 76.760 ;
        RECT 111.010 74.600 112.420 76.760 ;
        RECT 112.630 74.600 114.040 76.760 ;
        RECT 114.250 74.600 115.660 76.760 ;
        RECT 115.870 74.600 117.280 76.760 ;
        RECT 117.490 74.600 118.900 76.760 ;
        RECT 119.240 75.000 121.400 76.410 ;
        RECT 126.840 75.000 129.000 76.410 ;
        RECT 75.015 74.120 91.025 74.290 ;
        RECT 52.710 72.590 53.010 72.920 ;
        RECT 52.770 72.575 52.940 72.590 ;
        RECT 53.310 72.230 53.480 73.575 ;
        RECT 53.740 72.575 53.910 73.750 ;
        RECT 55.205 73.720 55.790 74.040 ;
        RECT 54.170 72.230 54.340 73.575 ;
        RECT 54.775 72.230 54.945 73.575 ;
        RECT 55.205 72.575 55.375 73.720 ;
        RECT 57.230 73.140 91.940 73.310 ;
        RECT 57.230 72.720 57.400 73.140 ;
        RECT 57.230 72.450 65.525 72.720 ;
        RECT 57.230 72.230 57.400 72.450 ;
        RECT 50.250 71.930 57.400 72.230 ;
        RECT 50.250 62.960 50.420 71.930 ;
        RECT 54.410 71.400 54.750 71.750 ;
        RECT 50.250 62.790 50.565 62.960 ;
        RECT 50.395 62.370 50.565 62.790 ;
        RECT 45.640 62.100 50.565 62.370 ;
        RECT 45.640 61.535 46.885 62.100 ;
        RECT 50.395 61.535 50.565 62.100 ;
        RECT 45.640 61.510 50.565 61.535 ;
        RECT 46.715 61.365 50.565 61.510 ;
        RECT 57.230 56.160 57.400 71.930 ;
        RECT 58.205 65.090 58.375 72.090 ;
        RECT 59.985 65.090 60.155 72.090 ;
        RECT 61.765 65.090 61.935 72.090 ;
        RECT 63.545 65.090 63.715 72.090 ;
        RECT 65.325 71.070 65.495 72.090 ;
        RECT 65.325 70.770 65.750 71.070 ;
        RECT 65.325 65.090 65.495 70.770 ;
        RECT 66.270 66.050 66.440 73.140 ;
        RECT 66.710 72.800 66.880 73.140 ;
        RECT 91.770 72.800 91.940 73.140 ;
        RECT 66.690 72.570 70.035 72.800 ;
        RECT 70.315 72.570 72.815 72.800 ;
        RECT 73.095 72.570 75.595 72.800 ;
        RECT 76.180 72.570 78.905 72.800 ;
        RECT 79.185 72.570 82.015 72.800 ;
        RECT 82.485 72.570 84.985 72.800 ;
        RECT 85.795 72.570 88.295 72.800 ;
        RECT 88.575 72.570 91.940 72.800 ;
        RECT 66.710 66.730 66.880 72.570 ;
        RECT 67.310 66.730 67.480 72.570 ;
        RECT 70.090 66.730 70.260 72.360 ;
        RECT 72.870 67.090 73.040 72.360 ;
        RECT 75.650 66.730 75.820 72.360 ;
        RECT 76.180 67.090 76.350 72.570 ;
        RECT 78.960 66.730 79.130 72.360 ;
        RECT 81.740 67.090 81.910 72.570 ;
        RECT 82.260 66.730 82.430 72.360 ;
        RECT 85.040 67.090 85.210 72.360 ;
        RECT 85.570 67.090 85.740 72.360 ;
        RECT 88.350 66.730 88.520 72.360 ;
        RECT 91.130 66.730 91.300 72.570 ;
        RECT 91.770 66.730 91.940 72.570 ;
        RECT 92.520 72.390 93.930 74.550 ;
        RECT 94.140 72.390 95.550 74.550 ;
        RECT 95.760 72.390 97.170 74.550 ;
        RECT 97.390 72.260 98.800 74.420 ;
        RECT 99.010 72.260 100.420 74.420 ;
        RECT 100.630 72.260 102.040 74.420 ;
        RECT 102.250 72.260 103.660 74.420 ;
        RECT 103.870 72.260 105.280 74.420 ;
        RECT 119.240 73.350 121.400 74.760 ;
        RECT 126.840 73.350 129.000 74.760 ;
        RECT 92.530 69.840 93.940 72.000 ;
        RECT 94.150 69.840 95.560 72.000 ;
        RECT 95.770 69.840 97.180 72.000 ;
        RECT 97.390 69.840 98.800 72.000 ;
        RECT 99.010 69.840 100.420 72.000 ;
        RECT 100.630 69.840 102.040 72.000 ;
        RECT 102.250 69.840 103.660 72.000 ;
        RECT 103.870 69.840 105.280 72.000 ;
        RECT 106.150 70.240 107.560 72.400 ;
        RECT 107.770 70.240 109.180 72.400 ;
        RECT 109.390 70.240 110.800 72.400 ;
        RECT 111.010 70.240 112.420 72.400 ;
        RECT 112.630 70.240 114.040 72.400 ;
        RECT 114.250 70.240 115.660 72.400 ;
        RECT 115.870 70.240 117.280 72.400 ;
        RECT 117.490 70.240 118.900 72.400 ;
        RECT 119.240 71.700 121.400 73.110 ;
        RECT 126.840 71.700 129.000 73.110 ;
        RECT 119.240 70.040 121.400 71.450 ;
        RECT 126.840 70.040 129.000 71.450 ;
        RECT 119.240 68.400 121.400 69.810 ;
        RECT 126.840 68.400 129.000 69.810 ;
        RECT 66.710 66.460 91.940 66.730 ;
        RECT 66.710 66.050 66.880 66.460 ;
        RECT 73.400 66.050 83.340 66.060 ;
        RECT 91.770 66.050 91.940 66.460 ;
        RECT 66.270 65.880 91.940 66.050 ;
        RECT 58.430 64.650 59.930 64.880 ;
        RECT 60.210 64.650 61.710 64.880 ;
        RECT 61.990 64.650 63.490 64.880 ;
        RECT 63.770 64.650 65.270 64.880 ;
        RECT 58.430 63.730 59.930 63.960 ;
        RECT 60.210 63.730 61.710 63.960 ;
        RECT 61.990 63.730 63.490 63.960 ;
        RECT 63.770 63.730 65.270 63.960 ;
        RECT 58.205 56.520 58.375 63.520 ;
        RECT 59.985 58.890 60.155 63.520 ;
        RECT 59.980 57.120 60.160 58.890 ;
        RECT 59.985 56.520 60.155 57.120 ;
        RECT 61.765 56.520 61.935 63.520 ;
        RECT 63.545 56.520 63.715 63.520 ;
        RECT 65.325 56.520 65.495 63.520 ;
        RECT 66.270 56.160 66.440 65.880 ;
        RECT 67.670 64.605 68.670 65.880 ;
        RECT 73.400 64.860 83.340 65.880 ;
        RECT 92.530 65.150 93.940 67.310 ;
        RECT 94.150 65.150 95.560 67.310 ;
        RECT 95.770 65.150 97.180 67.310 ;
        RECT 97.390 65.150 98.800 67.310 ;
        RECT 99.010 65.150 100.420 67.310 ;
        RECT 100.630 65.150 102.040 67.310 ;
        RECT 102.250 65.150 103.660 67.310 ;
        RECT 103.870 65.150 105.280 67.310 ;
        RECT 119.240 66.750 121.400 68.160 ;
        RECT 126.840 66.750 129.000 68.160 ;
        RECT 119.240 65.100 121.400 66.510 ;
        RECT 126.840 65.100 129.000 66.510 ;
        RECT 73.400 64.850 83.160 64.860 ;
        RECT 66.940 63.810 67.290 64.150 ;
        RECT 67.670 64.115 69.560 64.285 ;
        RECT 67.670 63.685 68.670 63.855 ;
        RECT 73.400 63.540 73.570 64.850 ;
        RECT 74.050 64.020 76.210 64.370 ;
        RECT 80.350 64.020 82.510 64.370 ;
        RECT 82.990 63.540 83.160 64.850 ;
        RECT 73.400 63.370 83.160 63.540 ;
        RECT 119.240 63.450 121.400 64.860 ;
        RECT 126.840 63.450 129.000 64.860 ;
        RECT 67.490 60.560 68.900 62.720 ;
        RECT 69.140 60.560 70.550 62.720 ;
        RECT 75.040 60.560 76.450 62.720 ;
        RECT 76.690 60.560 78.100 62.720 ;
        RECT 57.230 55.890 66.440 56.160 ;
        RECT 57.230 55.470 57.400 55.890 ;
        RECT 66.270 55.470 66.440 55.890 ;
        RECT 57.230 55.300 66.440 55.470 ;
        RECT 57.230 51.000 58.260 55.300 ;
        RECT 71.240 52.490 74.350 54.650 ;
        RECT 45.970 50.505 65.290 51.000 ;
        RECT 45.970 45.055 46.465 50.505 ;
        RECT 46.785 49.825 51.595 50.185 ;
        RECT 46.785 45.735 47.145 49.825 ;
        RECT 47.455 46.045 50.925 49.515 ;
        RECT 51.235 45.735 51.595 49.825 ;
        RECT 46.785 45.375 51.595 45.735 ;
        RECT 51.240 45.055 51.590 45.375 ;
        RECT 51.915 45.055 52.905 50.505 ;
        RECT 53.225 49.825 58.035 50.185 ;
        RECT 53.225 45.735 53.585 49.825 ;
        RECT 53.895 46.045 57.365 49.515 ;
        RECT 57.675 45.735 58.035 49.825 ;
        RECT 53.225 45.375 58.035 45.735 ;
        RECT 53.230 45.055 53.580 45.375 ;
        RECT 57.680 45.055 58.030 45.375 ;
        RECT 58.355 45.055 59.345 50.505 ;
        RECT 59.665 49.825 64.475 50.185 ;
        RECT 59.665 45.735 60.025 49.825 ;
        RECT 60.335 46.045 63.805 49.515 ;
        RECT 64.115 46.060 64.475 49.825 ;
        RECT 64.115 45.735 64.480 46.060 ;
        RECT 59.665 45.375 64.480 45.735 ;
        RECT 59.670 45.055 60.020 45.375 ;
        RECT 64.130 45.055 64.480 45.375 ;
        RECT 64.795 45.055 65.290 50.505 ;
        RECT 71.240 45.290 72.650 50.360 ;
        RECT 72.940 48.200 74.350 50.360 ;
        RECT 72.940 45.290 74.350 47.450 ;
        RECT 45.970 44.065 65.290 45.055 ;
        RECT 45.970 38.615 46.465 44.065 ;
        RECT 51.240 43.745 51.590 44.065 ;
        RECT 46.785 43.385 51.595 43.745 ;
        RECT 46.785 39.295 47.145 43.385 ;
        RECT 47.455 39.605 50.925 43.075 ;
        RECT 51.235 39.295 51.595 43.385 ;
        RECT 46.785 38.935 51.595 39.295 ;
        RECT 51.240 38.615 51.590 38.935 ;
        RECT 51.915 38.615 52.905 44.065 ;
        RECT 53.230 43.745 53.580 44.065 ;
        RECT 57.680 43.745 58.030 44.065 ;
        RECT 53.225 43.385 58.035 43.745 ;
        RECT 53.225 39.295 53.585 43.385 ;
        RECT 53.895 39.605 57.365 43.075 ;
        RECT 57.675 39.295 58.035 43.385 ;
        RECT 53.225 38.935 58.035 39.295 ;
        RECT 53.230 38.615 53.580 38.935 ;
        RECT 57.680 38.615 58.030 38.935 ;
        RECT 58.355 38.615 59.345 44.065 ;
        RECT 59.670 43.745 60.020 44.065 ;
        RECT 64.130 43.745 64.480 44.065 ;
        RECT 59.665 43.385 64.480 43.745 ;
        RECT 59.665 39.295 60.025 43.385 ;
        RECT 60.335 39.605 63.805 43.075 ;
        RECT 64.115 39.295 64.480 43.385 ;
        RECT 59.665 38.935 64.480 39.295 ;
        RECT 59.670 38.615 60.020 38.935 ;
        RECT 64.130 38.615 64.480 38.935 ;
        RECT 64.795 38.615 65.290 44.065 ;
        RECT 71.240 41.000 74.350 43.160 ;
        RECT 45.970 37.625 65.290 38.615 ;
        RECT 45.970 32.175 46.465 37.625 ;
        RECT 51.240 37.305 51.590 37.625 ;
        RECT 46.785 36.945 51.595 37.305 ;
        RECT 46.785 32.855 47.145 36.945 ;
        RECT 47.455 33.165 50.925 36.635 ;
        RECT 51.235 32.855 51.595 36.945 ;
        RECT 46.785 32.495 51.595 32.855 ;
        RECT 51.915 32.175 52.905 37.625 ;
        RECT 53.230 37.305 53.580 37.625 ;
        RECT 57.680 37.305 58.030 37.625 ;
        RECT 53.225 36.945 58.035 37.305 ;
        RECT 53.225 32.855 53.585 36.945 ;
        RECT 53.895 33.165 57.365 36.635 ;
        RECT 57.675 32.855 58.035 36.945 ;
        RECT 53.225 32.495 58.035 32.855 ;
        RECT 58.355 32.175 59.345 37.625 ;
        RECT 59.670 37.305 60.020 37.625 ;
        RECT 64.130 37.305 64.480 37.625 ;
        RECT 59.665 36.950 64.480 37.305 ;
        RECT 59.665 36.945 64.475 36.950 ;
        RECT 59.665 32.855 60.025 36.945 ;
        RECT 60.335 33.165 63.805 36.635 ;
        RECT 64.115 32.855 64.475 36.945 ;
        RECT 59.665 32.495 64.475 32.855 ;
        RECT 64.795 36.020 65.290 37.625 ;
        RECT 67.490 37.450 68.900 39.610 ;
        RECT 69.140 37.450 70.550 39.610 ;
        RECT 75.040 37.450 76.450 39.610 ;
        RECT 76.690 37.450 78.100 39.610 ;
        RECT 64.795 33.860 68.900 36.020 ;
        RECT 69.140 33.860 70.550 36.020 ;
        RECT 75.040 33.860 76.450 36.020 ;
        RECT 64.795 32.180 65.290 33.860 ;
        RECT 76.690 32.180 78.100 36.020 ;
        RECT 64.680 32.175 78.100 32.180 ;
        RECT 45.970 31.680 78.100 32.175 ;
        RECT 67.490 10.750 68.900 12.910 ;
        RECT 69.140 10.750 70.550 12.910 ;
        RECT 75.040 10.750 76.450 12.910 ;
        RECT 76.690 10.750 78.100 12.910 ;
      LAYER met1 ;
        RECT 47.855 187.460 76.440 187.550 ;
        RECT 47.855 187.280 118.595 187.460 ;
        RECT 76.170 187.190 118.595 187.280 ;
        RECT 92.125 187.180 92.395 187.190 ;
        RECT 54.950 181.870 68.290 182.880 ;
        RECT 28.070 180.100 28.320 180.890 ;
        RECT 28.030 179.530 28.380 180.100 ;
        RECT 28.070 178.785 28.320 179.530 ;
        RECT 28.610 178.790 29.460 180.900 ;
        RECT 28.630 178.785 28.880 178.790 ;
        RECT 29.190 178.785 29.440 178.790 ;
        RECT 29.720 178.780 30.570 180.890 ;
        RECT 30.850 178.780 31.700 180.890 ;
        RECT 31.970 178.780 32.820 180.890 ;
        RECT 33.110 180.100 33.360 180.890 ;
        RECT 33.110 179.500 36.210 180.100 ;
        RECT 37.880 179.530 38.380 180.100 ;
        RECT 33.110 178.785 33.360 179.500 ;
        RECT 35.710 178.830 36.210 179.500 ;
        RECT 37.260 172.535 37.810 172.980 ;
        RECT 35.710 167.685 36.710 167.955 ;
        RECT 35.250 165.900 35.520 167.230 ;
        RECT 38.000 166.990 38.270 179.530 ;
        RECT 51.135 179.490 72.105 180.500 ;
        RECT 76.985 179.820 77.355 180.080 ;
        RECT 80.305 180.035 80.595 180.065 ;
        RECT 86.865 180.035 87.155 180.065 ;
        RECT 80.305 179.865 87.155 180.035 ;
        RECT 80.305 179.835 80.595 179.865 ;
        RECT 86.865 179.835 87.155 179.865 ;
        RECT 90.130 179.820 90.450 180.080 ;
        RECT 92.110 179.775 92.370 180.145 ;
        RECT 95.375 179.810 102.195 180.100 ;
        RECT 105.200 179.830 105.520 180.090 ;
        RECT 118.320 179.830 118.640 180.090 ;
        RECT 47.840 176.285 48.100 176.605 ;
        RECT 75.140 176.285 75.400 176.605 ;
        RECT 71.330 175.060 71.590 175.075 ;
        RECT 51.660 174.735 51.920 175.060 ;
        RECT 71.320 174.755 71.590 175.060 ;
        RECT 71.320 174.740 71.580 174.755 ;
        RECT 90.160 173.020 90.420 173.670 ;
        RECT 118.350 173.040 118.610 176.570 ;
        RECT 38.460 172.535 39.010 172.980 ;
        RECT 48.110 172.610 54.920 172.880 ;
        RECT 55.200 172.610 68.040 172.880 ;
        RECT 68.320 172.610 80.310 172.880 ;
        RECT 80.590 172.610 86.870 172.880 ;
        RECT 87.150 172.610 95.380 172.880 ;
        RECT 95.660 172.610 101.940 172.880 ;
        RECT 102.220 172.610 105.220 172.880 ;
        RECT 105.500 172.610 118.340 172.880 ;
        RECT 45.070 171.590 46.760 172.240 ;
        RECT 61.780 171.405 62.790 172.610 ;
        RECT 83.605 172.045 83.875 172.610 ;
        RECT 87.450 171.870 87.850 172.610 ;
        RECT 98.670 172.045 98.940 172.610 ;
        RECT 82.500 171.670 87.850 171.870 ;
        RECT 59.785 170.970 63.855 171.240 ;
        RECT 48.285 170.685 57.845 170.955 ;
        RECT 65.455 170.880 80.025 171.150 ;
        RECT 42.915 167.955 43.295 168.315 ;
        RECT 44.320 167.735 44.640 167.760 ;
        RECT 39.400 167.465 45.345 167.735 ;
        RECT 44.320 167.440 44.640 167.465 ;
        RECT 48.285 167.305 48.555 170.685 ;
        RECT 53.200 167.500 53.460 168.780 ;
        RECT 57.575 167.305 57.845 170.685 ;
        RECT 61.780 169.515 62.790 170.630 ;
        RECT 61.065 168.505 63.855 169.515 ;
        RECT 69.330 167.955 69.590 170.515 ;
        RECT 82.500 169.400 83.810 171.670 ;
        RECT 75.140 168.540 83.810 169.400 ;
        RECT 84.070 169.290 87.100 171.450 ;
        RECT 87.310 169.290 90.340 171.450 ;
        RECT 90.550 169.290 93.580 171.450 ;
        RECT 93.840 170.970 95.150 171.430 ;
        RECT 96.700 171.295 96.960 171.615 ;
        RECT 93.840 169.960 96.220 170.970 ;
        RECT 106.865 170.965 107.135 172.610 ;
        RECT 96.735 169.965 107.135 170.965 ;
        RECT 93.840 169.325 95.150 169.960 ;
        RECT 96.680 168.610 96.970 169.480 ;
        RECT 48.285 167.035 51.380 167.305 ;
        RECT 51.660 167.035 54.470 167.305 ;
        RECT 54.750 167.035 57.845 167.305 ;
        RECT 38.460 166.940 39.010 166.965 ;
        RECT 40.170 166.940 40.470 167.030 ;
        RECT 75.140 166.965 75.860 168.540 ;
        RECT 38.460 166.760 40.470 166.940 ;
        RECT 37.490 165.940 37.920 165.990 ;
        RECT 37.490 165.900 37.950 165.940 ;
        RECT 35.250 165.640 37.950 165.900 ;
        RECT 28.060 159.290 28.910 161.400 ;
        RECT 29.190 161.390 29.440 161.395 ;
        RECT 29.750 161.390 30.000 161.395 ;
        RECT 29.180 159.280 30.030 161.390 ;
        RECT 30.290 159.290 31.120 161.400 ;
        RECT 31.410 159.290 32.260 161.400 ;
        RECT 32.540 159.290 33.390 161.400 ;
        RECT 35.250 159.615 35.520 165.640 ;
        RECT 37.490 165.600 37.950 165.640 ;
        RECT 37.490 165.580 37.920 165.600 ;
        RECT 38.460 165.465 39.010 166.760 ;
        RECT 40.170 166.700 40.470 166.760 ;
        RECT 60.040 166.610 63.600 166.880 ;
        RECT 65.710 166.695 68.710 166.965 ;
        RECT 69.600 166.695 75.880 166.965 ;
        RECT 76.770 166.695 79.770 166.965 ;
        RECT 46.280 165.920 46.780 166.130 ;
        RECT 45.310 165.600 46.780 165.920 ;
        RECT 35.775 164.625 36.145 164.885 ;
        RECT 36.830 164.670 37.230 165.120 ;
        RECT 38.460 164.955 39.505 165.465 ;
        RECT 46.280 165.450 46.780 165.600 ;
        RECT 38.460 164.820 39.180 164.955 ;
        RECT 42.640 164.460 42.960 164.810 ;
        RECT 78.995 164.700 79.550 164.720 ;
        RECT 56.370 164.600 59.975 164.700 ;
        RECT 48.115 164.430 59.975 164.600 ;
        RECT 60.190 164.430 78.235 164.700 ;
        RECT 78.515 164.680 81.015 164.700 ;
        RECT 78.515 164.450 81.880 164.680 ;
        RECT 78.515 164.430 81.015 164.450 ;
        RECT 48.115 164.330 56.640 164.430 ;
        RECT 43.690 164.095 44.000 164.100 ;
        RECT 45.250 164.095 47.010 164.100 ;
        RECT 40.780 163.825 41.800 164.095 ;
        RECT 42.250 163.825 42.910 164.095 ;
        RECT 43.220 163.825 44.310 164.095 ;
        RECT 44.685 163.825 47.010 164.095 ;
        RECT 43.670 163.820 44.130 163.825 ;
        RECT 45.250 163.820 47.010 163.825 ;
        RECT 47.550 163.685 47.810 164.005 ;
        RECT 44.350 163.280 44.690 163.630 ;
        RECT 47.610 159.190 47.750 163.685 ;
        RECT 55.350 162.650 55.700 162.950 ;
        RECT 74.935 162.640 75.195 162.960 ;
        RECT 82.500 162.260 83.810 166.745 ;
        RECT 84.120 162.265 85.430 166.745 ;
        RECT 85.740 162.265 87.050 166.745 ;
        RECT 87.360 162.265 88.670 166.745 ;
        RECT 88.980 162.260 90.290 166.745 ;
        RECT 90.600 162.265 91.910 166.745 ;
        RECT 92.220 162.260 93.530 166.745 ;
        RECT 93.840 162.265 95.150 166.745 ;
        RECT 96.140 166.505 97.450 168.610 ;
        RECT 97.760 166.500 100.690 168.610 ;
        RECT 101.000 166.500 103.930 168.610 ;
        RECT 104.240 166.500 107.170 168.610 ;
        RECT 107.480 166.505 108.790 168.610 ;
        RECT 109.180 165.230 111.340 168.290 ;
        RECT 116.805 166.930 118.910 168.240 ;
        RECT 96.140 164.250 97.450 164.255 ;
        RECT 97.760 164.250 99.070 164.255 ;
        RECT 96.140 162.140 99.070 164.250 ;
        RECT 99.380 162.150 102.310 164.260 ;
        RECT 102.620 162.150 105.550 164.260 ;
        RECT 105.860 164.255 107.480 164.260 ;
        RECT 105.860 162.150 108.790 164.255 ;
        RECT 55.790 161.730 56.050 162.050 ;
        RECT 109.180 161.920 111.340 164.980 ;
        RECT 116.780 163.580 118.940 166.640 ;
        RECT 49.895 159.980 50.125 160.055 ;
        RECT 55.840 159.980 55.980 161.730 ;
        RECT 62.765 161.425 63.025 161.795 ;
        RECT 75.435 161.480 75.755 161.740 ;
        RECT 49.895 159.840 55.980 159.980 ;
        RECT 49.895 159.765 50.125 159.840 ;
        RECT 53.455 159.190 53.685 159.265 ;
        RECT 35.710 158.560 37.620 159.070 ;
        RECT 47.610 159.050 53.685 159.190 ;
        RECT 33.310 154.250 36.830 154.610 ;
        RECT 33.310 153.980 39.770 154.250 ;
        RECT 33.310 153.430 36.830 153.980 ;
        RECT 33.310 153.420 36.820 153.430 ;
        RECT 47.610 152.530 47.750 159.050 ;
        RECT 53.455 158.975 53.685 159.050 ;
        RECT 48.115 157.410 55.575 158.420 ;
        RECT 48.345 156.510 51.650 156.780 ;
        RECT 51.930 156.510 55.235 156.780 ;
        RECT 53.435 156.325 53.705 156.510 ;
        RECT 49.870 156.055 53.705 156.325 ;
        RECT 49.870 155.860 50.140 156.055 ;
        RECT 48.370 155.590 51.650 155.860 ;
        RECT 51.930 155.590 55.210 155.860 ;
        RECT 55.435 154.960 55.575 157.410 ;
        RECT 47.975 153.950 55.575 154.960 ;
        RECT 53.455 153.300 53.685 153.375 ;
        RECT 55.840 153.300 55.980 159.840 ;
        RECT 80.910 158.610 81.270 158.660 ;
        RECT 57.220 158.340 81.270 158.610 ;
        RECT 80.910 158.310 81.270 158.340 ;
        RECT 82.500 157.580 85.440 159.690 ;
        RECT 85.740 157.580 88.680 159.690 ;
        RECT 88.970 157.580 91.910 159.690 ;
        RECT 92.220 157.580 95.160 159.690 ;
        RECT 109.180 158.630 111.340 161.690 ;
        RECT 116.780 160.280 118.940 163.340 ;
        RECT 57.610 156.485 58.610 156.755 ;
        RECT 82.150 156.250 84.320 156.780 ;
        RECT 56.880 155.690 57.230 156.030 ;
        RECT 59.270 155.900 66.150 156.250 ;
        RECT 70.290 155.900 84.320 156.250 ;
        RECT 57.795 155.740 58.475 155.765 ;
        RECT 57.610 155.330 58.610 155.740 ;
        RECT 82.150 155.360 84.320 155.900 ;
        RECT 109.180 155.330 111.340 158.390 ;
        RECT 116.780 156.980 118.940 160.040 ;
        RECT 116.805 155.380 118.910 156.690 ;
        RECT 53.455 153.160 55.980 153.300 ;
        RECT 53.455 153.085 53.685 153.160 ;
        RECT 49.895 152.530 50.125 152.605 ;
        RECT 47.610 152.390 50.125 152.530 ;
        RECT 57.430 152.440 60.490 154.600 ;
        RECT 64.980 152.440 68.040 154.600 ;
        RECT 49.895 152.315 50.125 152.390 ;
        RECT 49.870 151.000 50.150 151.010 ;
        RECT 49.870 148.920 50.240 151.000 ;
        RECT 48.115 147.770 55.465 148.040 ;
        RECT 48.345 146.920 58.810 147.190 ;
        RECT 37.600 138.100 53.540 141.190 ;
        RECT 37.600 128.340 40.660 138.100 ;
        RECT 44.045 131.695 47.095 134.745 ;
        RECT 50.480 128.340 53.540 138.100 ;
        RECT 57.480 137.710 58.810 146.920 ;
        RECT 61.230 144.395 62.540 146.500 ;
        RECT 62.930 144.395 64.240 146.500 ;
        RECT 61.230 140.110 62.540 142.215 ;
        RECT 62.930 140.110 67.990 142.240 ;
        RECT 57.480 129.360 58.790 137.710 ;
        RECT 61.230 137.195 62.540 139.300 ;
        RECT 62.930 137.195 64.240 139.300 ;
        RECT 61.230 132.910 62.540 135.015 ;
        RECT 62.930 132.910 64.240 135.015 ;
        RECT 59.130 129.360 60.440 131.465 ;
        RECT 65.030 129.360 66.340 131.465 ;
        RECT 66.680 129.360 67.990 140.110 ;
        RECT 65.030 128.980 66.330 129.360 ;
        RECT 37.600 125.250 54.170 128.340 ;
        RECT 59.130 128.180 66.330 128.980 ;
        RECT 57.480 125.765 58.790 127.870 ;
        RECT 59.130 125.765 60.440 128.180 ;
        RECT 65.030 125.765 66.340 127.870 ;
        RECT 66.680 125.765 67.990 127.870 ;
        RECT 57.430 102.630 60.490 104.790 ;
        RECT 64.980 102.630 68.040 104.790 ;
        RECT 57.915 95.580 86.500 95.670 ;
        RECT 128.540 95.580 129.010 95.600 ;
        RECT 57.915 95.400 129.010 95.580 ;
        RECT 86.230 95.310 129.010 95.400 ;
        RECT 102.185 95.300 102.455 95.310 ;
        RECT 128.540 95.290 129.010 95.310 ;
        RECT 65.010 89.990 78.350 91.000 ;
        RECT 38.130 88.220 38.380 89.010 ;
        RECT 38.090 87.650 38.440 88.220 ;
        RECT 38.130 86.905 38.380 87.650 ;
        RECT 38.670 86.910 39.520 89.020 ;
        RECT 38.690 86.905 38.940 86.910 ;
        RECT 39.250 86.905 39.500 86.910 ;
        RECT 39.780 86.900 40.630 89.010 ;
        RECT 40.910 86.900 41.760 89.010 ;
        RECT 42.030 86.900 42.880 89.010 ;
        RECT 43.170 88.220 43.420 89.010 ;
        RECT 43.170 87.620 46.270 88.220 ;
        RECT 47.940 87.650 48.440 88.220 ;
        RECT 43.170 86.905 43.420 87.620 ;
        RECT 45.770 86.950 46.270 87.620 ;
        RECT 47.320 80.655 47.870 81.100 ;
        RECT 45.770 75.805 46.770 76.075 ;
        RECT 45.310 74.020 45.580 75.350 ;
        RECT 48.060 75.110 48.330 87.650 ;
        RECT 61.195 87.610 82.165 88.620 ;
        RECT 87.045 87.940 87.415 88.200 ;
        RECT 90.365 88.155 90.655 88.185 ;
        RECT 96.925 88.155 97.215 88.185 ;
        RECT 90.365 87.985 97.215 88.155 ;
        RECT 90.365 87.955 90.655 87.985 ;
        RECT 96.925 87.955 97.215 87.985 ;
        RECT 100.190 87.940 100.510 88.200 ;
        RECT 102.170 87.895 102.430 88.265 ;
        RECT 105.435 87.930 112.255 88.220 ;
        RECT 115.260 87.950 115.580 88.210 ;
        RECT 128.380 87.950 128.700 88.210 ;
        RECT 57.900 84.405 58.160 84.725 ;
        RECT 85.200 84.405 85.460 84.725 ;
        RECT 81.390 83.180 81.650 83.195 ;
        RECT 61.720 82.855 61.980 83.180 ;
        RECT 81.380 82.875 81.650 83.180 ;
        RECT 81.380 82.860 81.640 82.875 ;
        RECT 100.220 81.140 100.480 81.790 ;
        RECT 128.410 81.160 128.670 84.690 ;
        RECT 48.520 80.655 49.070 81.100 ;
        RECT 58.170 80.730 64.980 81.000 ;
        RECT 65.260 80.730 78.100 81.000 ;
        RECT 78.380 80.730 90.370 81.000 ;
        RECT 90.650 80.730 96.930 81.000 ;
        RECT 97.210 80.730 105.440 81.000 ;
        RECT 105.720 80.730 112.000 81.000 ;
        RECT 112.280 80.730 115.280 81.000 ;
        RECT 115.560 80.730 128.400 81.000 ;
        RECT 71.840 79.525 72.850 80.730 ;
        RECT 93.665 80.165 93.935 80.730 ;
        RECT 97.510 79.990 97.910 80.730 ;
        RECT 108.730 80.165 109.000 80.730 ;
        RECT 92.570 79.860 97.910 79.990 ;
        RECT 92.560 79.790 97.910 79.860 ;
        RECT 69.845 79.090 73.915 79.360 ;
        RECT 58.345 78.805 67.905 79.075 ;
        RECT 75.515 79.000 90.085 79.270 ;
        RECT 92.560 79.190 93.890 79.790 ;
        RECT 106.760 79.415 107.020 79.735 ;
        RECT 52.975 76.075 53.355 76.435 ;
        RECT 54.410 75.855 54.730 75.880 ;
        RECT 49.460 75.585 55.405 75.855 ;
        RECT 54.410 75.560 54.730 75.585 ;
        RECT 58.345 75.425 58.615 78.805 ;
        RECT 63.260 75.620 63.520 76.900 ;
        RECT 67.635 75.425 67.905 78.805 ;
        RECT 92.570 78.960 93.890 79.190 ;
        RECT 94.190 79.100 95.500 79.210 ;
        RECT 95.810 79.100 97.120 79.210 ;
        RECT 71.840 77.635 72.850 78.750 ;
        RECT 71.125 76.625 73.915 77.635 ;
        RECT 79.390 76.075 79.650 78.635 ;
        RECT 92.570 77.520 93.880 78.960 ;
        RECT 85.200 77.105 93.880 77.520 ;
        RECT 85.200 76.660 93.850 77.105 ;
        RECT 94.150 76.940 97.180 79.100 ;
        RECT 97.390 76.940 100.420 79.100 ;
        RECT 100.630 76.940 103.660 79.100 ;
        RECT 103.950 79.080 106.280 79.090 ;
        RECT 116.925 79.085 117.195 80.730 ;
        RECT 103.920 78.080 106.280 79.080 ;
        RECT 106.795 78.085 117.195 79.085 ;
        RECT 103.920 78.070 106.030 78.080 ;
        RECT 103.920 77.990 105.760 78.070 ;
        RECT 103.920 76.975 105.230 77.990 ;
        RECT 106.740 76.730 107.030 77.600 ;
        RECT 58.345 75.155 61.440 75.425 ;
        RECT 61.720 75.155 64.530 75.425 ;
        RECT 64.810 75.155 67.905 75.425 ;
        RECT 48.520 75.060 49.070 75.085 ;
        RECT 50.230 75.060 50.530 75.150 ;
        RECT 85.200 75.085 85.920 76.660 ;
        RECT 92.100 76.650 93.850 76.660 ;
        RECT 48.520 74.880 50.530 75.060 ;
        RECT 47.570 74.020 48.010 74.060 ;
        RECT 45.310 73.760 48.010 74.020 ;
        RECT 38.120 67.410 38.970 69.520 ;
        RECT 39.250 69.510 39.500 69.515 ;
        RECT 39.810 69.510 40.060 69.515 ;
        RECT 39.240 67.400 40.090 69.510 ;
        RECT 40.350 67.410 41.180 69.520 ;
        RECT 41.470 67.410 42.320 69.520 ;
        RECT 42.600 67.410 43.450 69.520 ;
        RECT 45.310 67.735 45.580 73.760 ;
        RECT 47.570 73.720 48.010 73.760 ;
        RECT 48.520 73.585 49.070 74.880 ;
        RECT 50.230 74.820 50.530 74.880 ;
        RECT 70.100 74.730 73.660 75.000 ;
        RECT 75.770 74.815 78.770 75.085 ;
        RECT 79.660 74.815 85.940 75.085 ;
        RECT 86.830 74.815 89.830 75.085 ;
        RECT 106.200 74.625 107.510 76.730 ;
        RECT 107.820 74.620 110.750 76.730 ;
        RECT 111.060 74.620 113.990 76.730 ;
        RECT 114.300 74.620 117.230 76.730 ;
        RECT 117.540 74.625 118.850 76.730 ;
        RECT 56.340 74.040 56.840 74.250 ;
        RECT 55.370 73.720 56.840 74.040 ;
        RECT 45.835 72.745 46.205 73.005 ;
        RECT 46.890 72.790 47.290 73.240 ;
        RECT 48.520 73.075 49.565 73.585 ;
        RECT 56.340 73.570 56.840 73.720 ;
        RECT 92.570 73.250 93.880 74.525 ;
        RECT 94.190 73.250 95.500 74.525 ;
        RECT 95.810 73.250 97.120 74.525 ;
        RECT 48.520 72.940 49.240 73.075 ;
        RECT 52.700 72.580 53.020 72.930 ;
        RECT 89.055 72.820 89.610 72.840 ;
        RECT 66.430 72.720 70.035 72.820 ;
        RECT 58.175 72.550 70.035 72.720 ;
        RECT 70.250 72.550 88.295 72.820 ;
        RECT 88.575 72.800 91.075 72.820 ;
        RECT 88.575 72.570 91.940 72.800 ;
        RECT 88.575 72.550 91.075 72.570 ;
        RECT 58.175 72.450 66.700 72.550 ;
        RECT 92.570 72.420 93.890 73.250 ;
        RECT 94.190 72.420 95.510 73.250 ;
        RECT 95.810 72.420 97.130 73.250 ;
        RECT 53.750 72.215 54.060 72.220 ;
        RECT 55.310 72.215 57.070 72.220 ;
        RECT 50.840 71.945 51.860 72.215 ;
        RECT 52.310 71.945 52.970 72.215 ;
        RECT 53.280 71.945 54.370 72.215 ;
        RECT 54.745 71.945 57.070 72.215 ;
        RECT 53.730 71.940 54.190 71.945 ;
        RECT 55.310 71.940 57.070 71.945 ;
        RECT 57.610 71.805 57.870 72.125 ;
        RECT 54.410 71.400 54.750 71.750 ;
        RECT 57.670 67.310 57.810 71.805 ;
        RECT 65.410 70.770 65.760 71.070 ;
        RECT 84.995 70.760 85.255 71.080 ;
        RECT 65.850 69.850 66.110 70.170 ;
        RECT 59.955 68.100 60.185 68.175 ;
        RECT 65.900 68.100 66.040 69.850 ;
        RECT 72.825 69.545 73.085 69.915 ;
        RECT 92.580 69.865 93.890 72.420 ;
        RECT 94.200 69.865 95.510 72.420 ;
        RECT 95.820 69.865 97.130 72.420 ;
        RECT 97.440 69.865 98.750 74.395 ;
        RECT 99.060 69.865 100.370 74.395 ;
        RECT 100.680 69.865 101.990 74.395 ;
        RECT 102.300 69.865 103.610 74.395 ;
        RECT 103.920 69.865 105.230 74.395 ;
        RECT 119.240 73.350 121.400 76.410 ;
        RECT 126.865 75.050 128.970 76.360 ;
        RECT 106.200 72.370 107.510 72.375 ;
        RECT 107.820 72.370 109.130 72.375 ;
        RECT 106.200 70.260 109.130 72.370 ;
        RECT 109.440 70.270 112.370 72.380 ;
        RECT 112.680 70.270 115.610 72.380 ;
        RECT 115.920 72.375 117.540 72.380 ;
        RECT 115.920 70.270 118.850 72.375 ;
        RECT 119.240 70.040 121.400 73.100 ;
        RECT 126.840 71.700 129.000 74.760 ;
        RECT 85.495 69.600 85.815 69.860 ;
        RECT 59.955 67.960 66.040 68.100 ;
        RECT 59.955 67.885 60.185 67.960 ;
        RECT 63.515 67.310 63.745 67.385 ;
        RECT 45.770 66.680 47.680 67.190 ;
        RECT 57.670 67.170 63.745 67.310 ;
        RECT 36.640 62.370 46.860 62.670 ;
        RECT 36.640 62.100 49.830 62.370 ;
        RECT 36.640 61.510 46.860 62.100 ;
        RECT 57.670 60.650 57.810 67.170 ;
        RECT 63.515 67.095 63.745 67.170 ;
        RECT 58.175 65.530 65.635 66.540 ;
        RECT 58.405 64.630 61.710 64.900 ;
        RECT 61.990 64.630 65.295 64.900 ;
        RECT 63.495 64.445 63.765 64.630 ;
        RECT 59.930 64.175 63.765 64.445 ;
        RECT 59.930 63.980 60.200 64.175 ;
        RECT 58.430 63.710 61.710 63.980 ;
        RECT 61.990 63.710 65.270 63.980 ;
        RECT 65.495 63.080 65.635 65.530 ;
        RECT 58.035 62.070 65.635 63.080 ;
        RECT 63.515 61.420 63.745 61.495 ;
        RECT 65.900 61.420 66.040 67.960 ;
        RECT 91.010 66.730 91.400 66.780 ;
        RECT 67.280 66.460 91.400 66.730 ;
        RECT 91.010 66.440 91.400 66.460 ;
        RECT 92.580 65.180 95.510 67.290 ;
        RECT 95.820 65.180 98.750 67.290 ;
        RECT 99.060 65.180 101.990 67.290 ;
        RECT 102.300 65.180 105.230 67.290 ;
        RECT 119.240 66.750 121.400 69.810 ;
        RECT 126.840 68.400 129.000 71.460 ;
        RECT 67.670 64.605 68.670 64.875 ;
        RECT 92.210 64.370 94.380 64.900 ;
        RECT 66.940 63.810 67.290 64.150 ;
        RECT 69.330 64.020 76.210 64.370 ;
        RECT 80.350 64.020 94.380 64.370 ;
        RECT 67.855 63.860 68.535 63.885 ;
        RECT 67.670 63.450 68.670 63.860 ;
        RECT 92.210 63.480 94.380 64.020 ;
        RECT 119.240 63.450 121.400 66.510 ;
        RECT 126.840 65.100 129.000 68.160 ;
        RECT 126.865 63.500 128.970 64.810 ;
        RECT 63.515 61.280 66.040 61.420 ;
        RECT 63.515 61.205 63.745 61.280 ;
        RECT 59.955 60.650 60.185 60.725 ;
        RECT 57.670 60.510 60.185 60.650 ;
        RECT 67.490 60.560 70.550 62.720 ;
        RECT 75.040 60.560 78.100 62.720 ;
        RECT 59.955 60.435 60.185 60.510 ;
        RECT 59.930 59.120 60.210 59.130 ;
        RECT 59.930 57.040 60.300 59.120 ;
        RECT 58.175 55.890 65.525 56.160 ;
        RECT 58.405 55.040 68.870 55.310 ;
        RECT 47.660 46.220 63.600 49.310 ;
        RECT 47.660 36.460 50.720 46.220 ;
        RECT 54.105 39.815 57.155 42.865 ;
        RECT 60.540 36.460 63.600 46.220 ;
        RECT 67.540 45.830 68.870 55.040 ;
        RECT 71.290 52.515 72.600 54.620 ;
        RECT 72.990 52.515 74.300 54.620 ;
        RECT 71.290 48.230 72.600 50.335 ;
        RECT 72.990 48.230 78.050 50.360 ;
        RECT 67.540 37.480 68.850 45.830 ;
        RECT 71.290 45.315 72.600 47.420 ;
        RECT 72.990 45.315 74.300 47.420 ;
        RECT 71.290 41.030 72.600 43.135 ;
        RECT 72.990 41.030 74.300 43.135 ;
        RECT 69.190 37.480 70.500 39.585 ;
        RECT 75.090 37.480 76.400 39.585 ;
        RECT 76.740 37.480 78.050 48.230 ;
        RECT 75.090 37.100 76.390 37.480 ;
        RECT 47.660 33.370 64.230 36.460 ;
        RECT 69.190 36.300 76.390 37.100 ;
        RECT 67.540 33.885 68.850 35.990 ;
        RECT 69.190 33.885 70.500 36.300 ;
        RECT 75.090 33.885 76.400 35.990 ;
        RECT 76.740 33.885 78.050 35.990 ;
        RECT 67.490 10.750 70.550 12.910 ;
        RECT 75.040 10.750 78.100 12.910 ;
      LAYER met2 ;
        RECT 27.980 179.530 38.380 180.100 ;
        RECT 77.010 180.035 77.330 180.080 ;
        RECT 90.130 180.035 90.450 180.080 ;
        RECT 77.010 179.865 90.450 180.035 ;
        RECT 77.010 179.820 77.330 179.865 ;
        RECT 90.130 179.820 90.450 179.865 ;
        RECT 92.080 180.045 92.400 180.090 ;
        RECT 105.200 180.045 105.520 180.090 ;
        RECT 118.320 180.045 118.640 180.090 ;
        RECT 92.080 179.875 118.640 180.045 ;
        RECT 92.080 179.830 92.400 179.875 ;
        RECT 105.200 179.830 105.520 179.875 ;
        RECT 118.320 179.830 118.640 179.875 ;
        RECT 35.710 164.610 36.210 179.230 ;
        RECT 47.830 176.260 48.110 176.630 ;
        RECT 75.130 176.260 75.410 176.630 ;
        RECT 118.350 176.380 118.610 176.405 ;
        RECT 51.645 174.710 51.930 175.080 ;
        RECT 71.320 175.060 71.600 175.100 ;
        RECT 71.320 174.730 71.625 175.060 ;
        RECT 71.345 174.690 71.625 174.730 ;
        RECT 90.150 173.025 90.430 173.665 ;
        RECT 53.545 172.610 69.750 172.880 ;
        RECT 78.940 172.610 88.535 172.880 ;
        RECT 93.730 172.610 103.955 172.880 ;
        RECT 45.030 171.560 45.510 172.280 ;
        RECT 61.780 172.070 98.965 172.340 ;
        RECT 61.780 169.730 62.790 172.070 ;
        RECT 42.840 167.880 43.360 168.390 ;
        RECT 44.240 167.350 44.720 167.840 ;
        RECT 53.200 167.810 53.460 168.780 ;
        RECT 47.610 167.670 60.585 167.810 ;
        RECT 37.430 165.520 37.950 166.020 ;
        RECT 46.280 165.450 46.780 166.130 ;
        RECT 36.830 164.670 37.230 165.120 ;
        RECT 42.640 164.460 42.960 164.810 ;
        RECT 42.670 163.630 42.930 164.460 ;
        RECT 47.610 164.005 47.750 167.670 ;
        RECT 53.200 167.500 53.460 167.670 ;
        RECT 53.490 167.235 54.450 167.295 ;
        RECT 55.780 167.235 55.980 167.240 ;
        RECT 53.490 167.095 55.980 167.235 ;
        RECT 53.490 167.035 54.450 167.095 ;
        RECT 55.700 167.090 55.980 167.095 ;
        RECT 48.365 165.400 48.645 165.770 ;
        RECT 54.935 165.410 55.215 165.780 ;
        RECT 47.550 163.685 47.810 164.005 ;
        RECT 42.670 163.280 44.690 163.630 ;
        RECT 33.300 153.420 34.880 154.610 ;
        RECT 48.370 146.895 48.640 165.400 ;
        RECT 49.870 156.325 50.140 156.805 ;
        RECT 49.870 156.055 53.745 156.325 ;
        RECT 53.475 155.565 53.745 156.055 ;
        RECT 49.870 148.920 50.240 151.010 ;
        RECT 54.940 147.480 55.210 165.410 ;
        RECT 55.350 162.620 55.670 163.000 ;
        RECT 55.840 162.050 55.980 167.090 ;
        RECT 60.445 166.905 60.585 167.670 ;
        RECT 60.385 166.585 60.645 166.905 ;
        RECT 55.790 161.730 56.050 162.050 ;
        RECT 62.735 161.695 63.055 169.460 ;
        RECT 69.330 167.955 69.590 170.515 ;
        RECT 93.830 168.560 95.150 171.420 ;
        RECT 96.690 171.270 96.970 171.640 ;
        RECT 69.375 164.695 69.545 167.955 ;
        RECT 93.830 166.430 108.790 168.560 ;
        RECT 117.780 168.290 118.610 176.380 ;
        RECT 116.780 166.880 118.940 168.290 ;
        RECT 66.840 164.435 71.475 164.695 ;
        RECT 74.925 162.615 75.205 162.985 ;
        RECT 75.435 161.695 75.755 161.740 ;
        RECT 62.735 161.525 75.755 161.695 ;
        RECT 62.735 156.250 63.055 161.525 ;
        RECT 75.435 161.480 75.755 161.525 ;
        RECT 107.480 158.700 108.790 166.430 ;
        RECT 80.850 158.250 108.790 158.700 ;
        RECT 56.860 155.670 57.250 156.050 ;
        RECT 62.730 155.900 63.060 156.250 ;
        RECT 57.610 155.330 58.610 155.740 ;
        RECT 82.150 155.360 84.320 156.780 ;
        RECT 107.480 156.690 108.790 158.250 ;
        RECT 107.480 155.380 118.910 156.690 ;
        RECT 54.940 147.180 64.250 147.480 ;
        RECT 57.610 144.580 58.610 145.260 ;
        RECT 62.930 140.110 64.250 147.180 ;
        RECT 51.470 137.190 64.240 139.300 ;
        RECT 44.930 132.550 58.790 133.780 ;
        RECT 57.480 129.350 58.790 132.550 ;
        RECT 59.130 129.360 60.440 131.460 ;
        RECT 59.130 128.980 60.430 129.360 ;
        RECT 59.130 128.180 66.330 128.980 ;
        RECT 65.030 127.870 66.330 128.180 ;
        RECT 65.030 125.770 66.340 127.870 ;
        RECT 128.580 95.210 129.060 95.670 ;
        RECT 38.040 87.650 48.440 88.220 ;
        RECT 87.070 88.155 87.390 88.200 ;
        RECT 100.190 88.155 100.510 88.200 ;
        RECT 87.070 87.985 100.510 88.155 ;
        RECT 87.070 87.940 87.390 87.985 ;
        RECT 100.190 87.940 100.510 87.985 ;
        RECT 102.140 88.165 102.460 88.210 ;
        RECT 115.260 88.165 115.580 88.210 ;
        RECT 128.380 88.165 128.700 88.210 ;
        RECT 102.140 87.995 128.700 88.165 ;
        RECT 102.140 87.950 102.460 87.995 ;
        RECT 115.260 87.950 115.580 87.995 ;
        RECT 128.380 87.950 128.700 87.995 ;
        RECT 45.770 72.730 46.270 87.350 ;
        RECT 57.890 84.380 58.170 84.750 ;
        RECT 85.190 84.380 85.470 84.750 ;
        RECT 128.410 84.500 128.670 84.525 ;
        RECT 61.705 82.830 61.990 83.200 ;
        RECT 81.380 83.180 81.660 83.220 ;
        RECT 81.380 82.850 81.685 83.180 ;
        RECT 81.405 82.810 81.685 82.850 ;
        RECT 100.210 81.145 100.490 81.785 ;
        RECT 63.605 80.730 79.810 81.000 ;
        RECT 89.000 80.730 98.595 81.000 ;
        RECT 103.790 80.730 114.015 81.000 ;
        RECT 71.840 80.190 109.025 80.460 ;
        RECT 71.840 77.850 72.850 80.190 ;
        RECT 106.750 79.390 107.030 79.760 ;
        RECT 52.950 76.030 53.380 76.480 ;
        RECT 54.310 75.460 54.830 75.980 ;
        RECT 63.260 75.930 63.520 76.900 ;
        RECT 57.670 75.790 70.645 75.930 ;
        RECT 47.500 73.650 47.990 74.130 ;
        RECT 56.340 73.570 56.840 74.250 ;
        RECT 46.890 72.790 47.290 73.240 ;
        RECT 52.700 72.580 53.020 72.930 ;
        RECT 52.730 71.750 52.990 72.580 ;
        RECT 57.670 72.125 57.810 75.790 ;
        RECT 63.260 75.620 63.520 75.790 ;
        RECT 63.550 75.355 64.510 75.415 ;
        RECT 65.840 75.355 66.040 75.360 ;
        RECT 63.550 75.215 66.040 75.355 ;
        RECT 63.550 75.155 64.510 75.215 ;
        RECT 65.760 75.210 66.040 75.215 ;
        RECT 58.425 73.520 58.705 73.890 ;
        RECT 64.995 73.530 65.275 73.900 ;
        RECT 57.610 71.805 57.870 72.125 ;
        RECT 52.730 71.400 54.750 71.750 ;
        RECT 36.870 61.650 37.760 62.540 ;
        RECT 58.430 55.015 58.700 73.520 ;
        RECT 59.930 64.445 60.200 64.925 ;
        RECT 59.930 64.175 63.805 64.445 ;
        RECT 63.535 63.685 63.805 64.175 ;
        RECT 59.930 57.040 60.300 59.130 ;
        RECT 65.000 55.600 65.270 73.530 ;
        RECT 65.410 70.740 65.730 71.120 ;
        RECT 65.900 70.170 66.040 75.210 ;
        RECT 70.505 75.025 70.645 75.790 ;
        RECT 70.445 74.705 70.705 75.025 ;
        RECT 65.850 69.850 66.110 70.170 ;
        RECT 72.795 69.815 73.115 77.580 ;
        RECT 79.390 76.075 79.650 78.635 ;
        RECT 103.910 76.680 105.230 79.070 ;
        RECT 79.435 72.815 79.605 76.075 ;
        RECT 103.910 74.550 118.850 76.680 ;
        RECT 127.840 76.410 128.670 84.500 ;
        RECT 126.840 75.000 129.000 76.410 ;
        RECT 76.900 72.555 81.535 72.815 ;
        RECT 84.985 70.735 85.265 71.105 ;
        RECT 85.495 69.815 85.815 69.860 ;
        RECT 72.795 69.645 85.815 69.815 ;
        RECT 72.795 64.370 73.115 69.645 ;
        RECT 85.495 69.600 85.815 69.645 ;
        RECT 117.540 66.780 118.850 74.550 ;
        RECT 91.010 66.440 118.850 66.780 ;
        RECT 66.920 63.790 67.310 64.170 ;
        RECT 72.790 64.020 73.120 64.370 ;
        RECT 67.670 63.450 68.670 63.860 ;
        RECT 92.210 63.480 94.380 64.900 ;
        RECT 117.540 64.810 118.850 66.440 ;
        RECT 117.540 63.500 128.970 64.810 ;
        RECT 65.000 55.300 74.310 55.600 ;
        RECT 67.670 52.700 68.670 53.380 ;
        RECT 72.990 48.230 74.310 55.300 ;
        RECT 61.530 45.310 74.300 47.420 ;
        RECT 54.990 40.670 68.850 41.900 ;
        RECT 67.540 37.470 68.850 40.670 ;
        RECT 69.190 37.480 70.500 39.580 ;
        RECT 69.190 37.100 70.490 37.480 ;
        RECT 69.190 36.300 76.390 37.100 ;
        RECT 75.090 35.990 76.390 36.300 ;
        RECT 75.090 33.890 76.400 35.990 ;
      LAYER met3 ;
        RECT 42.840 192.170 43.350 192.320 ;
        RECT 42.840 167.880 43.360 192.170 ;
        RECT 47.805 176.595 48.655 176.610 ;
        RECT 75.105 176.595 75.435 176.610 ;
        RECT 47.805 176.295 75.435 176.595 ;
        RECT 47.805 176.050 48.655 176.295 ;
        RECT 75.105 176.280 75.435 176.295 ;
        RECT 44.230 167.390 44.730 167.840 ;
        RECT 25.110 166.970 44.730 167.390 ;
        RECT 37.400 165.490 37.980 166.050 ;
        RECT 36.780 164.610 37.280 165.190 ;
        RECT 45.040 158.010 45.790 172.550 ;
        RECT 46.280 156.050 46.780 166.130 ;
        RECT 48.355 165.750 48.655 176.050 ;
        RECT 51.620 175.040 51.950 175.060 ;
        RECT 51.620 174.740 71.650 175.040 ;
        RECT 51.620 174.730 51.950 174.740 ;
        RECT 54.925 165.760 55.225 174.740 ;
        RECT 71.320 174.710 71.650 174.740 ;
        RECT 90.125 173.180 90.455 173.510 ;
        RECT 90.140 171.605 90.440 173.180 ;
        RECT 96.665 171.605 96.995 171.620 ;
        RECT 90.140 171.305 96.995 171.605 ;
        RECT 96.665 171.290 96.995 171.305 ;
        RECT 116.780 166.880 118.940 168.290 ;
        RECT 48.340 165.420 48.670 165.750 ;
        RECT 54.910 165.430 55.240 165.760 ;
        RECT 55.320 162.950 55.730 163.000 ;
        RECT 74.900 162.950 75.230 162.965 ;
        RECT 55.320 162.650 75.230 162.950 ;
        RECT 55.320 162.620 55.730 162.650 ;
        RECT 74.900 162.635 75.230 162.650 ;
        RECT 46.280 155.670 57.250 156.050 ;
        RECT 4.000 153.430 34.880 154.610 ;
        RECT 4.000 153.410 14.030 153.430 ;
        RECT 49.870 148.920 50.300 151.010 ;
        RECT 57.610 144.580 58.610 155.740 ;
        RECT 82.150 155.360 84.320 156.780 ;
        RECT 82.150 155.350 84.165 155.360 ;
        RECT 72.040 145.370 82.150 154.020 ;
        RECT 83.350 145.370 93.460 154.020 ;
        RECT 72.040 135.520 82.150 144.170 ;
        RECT 83.350 135.520 93.460 144.170 ;
        RECT 72.040 125.670 82.150 134.320 ;
        RECT 83.350 125.670 93.460 134.320 ;
        RECT 72.040 115.820 82.150 124.470 ;
        RECT 83.350 115.820 93.460 124.470 ;
        RECT 52.910 99.420 53.430 99.940 ;
        RECT 52.920 76.010 53.410 99.420 ;
        RECT 128.570 95.190 129.070 95.680 ;
        RECT 57.865 84.715 58.715 84.730 ;
        RECT 85.165 84.715 85.495 84.730 ;
        RECT 57.865 84.415 85.495 84.715 ;
        RECT 57.865 84.170 58.715 84.415 ;
        RECT 85.165 84.400 85.495 84.415 ;
        RECT 47.480 73.630 48.010 74.150 ;
        RECT 46.840 72.730 47.340 73.310 ;
        RECT 54.310 68.500 54.830 75.980 ;
        RECT 56.340 64.170 56.840 74.250 ;
        RECT 58.415 73.870 58.715 84.170 ;
        RECT 61.680 83.160 62.010 83.180 ;
        RECT 61.680 82.860 81.710 83.160 ;
        RECT 61.680 82.850 62.010 82.860 ;
        RECT 64.985 73.880 65.285 82.860 ;
        RECT 81.380 82.830 81.710 82.860 ;
        RECT 100.185 81.300 100.515 81.630 ;
        RECT 100.200 79.725 100.500 81.300 ;
        RECT 106.725 79.725 107.055 79.740 ;
        RECT 100.200 79.425 107.055 79.725 ;
        RECT 106.725 79.410 107.055 79.425 ;
        RECT 126.840 75.000 129.000 76.410 ;
        RECT 58.400 73.540 58.730 73.870 ;
        RECT 64.970 73.550 65.300 73.880 ;
        RECT 65.380 71.070 65.790 71.120 ;
        RECT 84.960 71.070 85.290 71.085 ;
        RECT 65.380 70.770 85.290 71.070 ;
        RECT 65.380 70.740 65.790 70.770 ;
        RECT 84.960 70.755 85.290 70.770 ;
        RECT 56.340 63.790 67.310 64.170 ;
        RECT 3.990 62.680 12.090 62.690 ;
        RECT 3.990 61.500 38.230 62.680 ;
        RECT 3.990 61.490 12.090 61.500 ;
        RECT 59.930 57.040 60.360 59.130 ;
        RECT 67.670 52.700 68.670 63.860 ;
        RECT 92.210 63.480 94.380 64.900 ;
        RECT 92.210 63.470 94.225 63.480 ;
        RECT 82.100 53.490 92.210 62.140 ;
        RECT 93.410 53.490 103.520 62.140 ;
        RECT 82.100 43.640 92.210 52.290 ;
        RECT 93.410 43.640 103.520 52.290 ;
        RECT 82.100 33.790 92.210 42.440 ;
        RECT 93.410 33.790 103.520 42.440 ;
        RECT 82.100 23.940 92.210 32.590 ;
        RECT 93.410 23.940 103.520 32.590 ;
      LAYER met4 ;
        RECT 56.705 219.525 57.205 220.025 ;
        RECT 56.705 219.025 57.705 219.525 ;
        RECT 58.605 219.485 59.175 220.045 ;
        RECT 58.075 219.025 59.175 219.485 ;
        RECT 56.705 218.525 59.175 219.025 ;
        RECT 56.705 216.525 57.205 218.525 ;
        RECT 57.705 218.485 59.175 218.525 ;
        RECT 57.705 218.025 58.205 218.485 ;
        RECT 58.605 216.545 59.175 218.485 ;
        RECT 59.565 219.635 62.005 220.065 ;
        RECT 59.565 218.625 60.135 219.635 ;
        RECT 61.435 218.625 62.005 219.635 ;
        RECT 59.565 218.195 62.005 218.625 ;
        RECT 59.565 216.565 60.135 218.195 ;
        RECT 61.435 216.565 62.005 218.195 ;
        RECT 63.055 219.525 63.555 220.025 ;
        RECT 63.055 219.025 64.055 219.525 ;
        RECT 64.955 219.485 65.525 220.045 ;
        RECT 64.425 219.025 65.525 219.485 ;
        RECT 63.055 218.525 65.525 219.025 ;
        RECT 63.055 216.525 63.555 218.525 ;
        RECT 64.055 218.485 65.525 218.525 ;
        RECT 64.055 218.025 64.555 218.485 ;
        RECT 64.955 216.545 65.525 218.485 ;
        RECT 65.855 219.635 68.075 220.065 ;
        RECT 65.855 218.555 66.425 219.635 ;
        RECT 68.675 219.525 70.675 220.025 ;
        RECT 65.855 218.125 68.065 218.555 ;
        RECT 65.855 216.995 66.425 218.125 ;
        RECT 68.675 217.025 69.175 219.525 ;
        RECT 70.175 219.025 71.175 219.525 ;
        RECT 70.675 217.525 71.175 219.025 ;
        RECT 70.175 217.025 71.175 217.525 ;
        RECT 71.645 218.485 72.145 219.985 ;
        RECT 73.145 218.485 73.645 219.985 ;
        RECT 71.645 217.985 73.645 218.485 ;
        RECT 65.845 216.565 68.055 216.995 ;
        RECT 68.675 216.525 70.675 217.025 ;
        RECT 71.645 216.485 72.145 217.985 ;
        RECT 73.145 216.485 73.645 217.985 ;
        RECT 74.145 219.565 76.585 219.995 ;
        RECT 74.145 218.555 74.715 219.565 ;
        RECT 76.015 218.555 76.585 219.565 ;
        RECT 74.145 218.125 76.585 218.555 ;
        RECT 74.145 216.495 74.715 218.125 ;
        RECT 76.015 216.495 76.585 218.125 ;
        RECT 46.605 210.415 47.605 214.415 ;
        RECT 51.105 213.415 54.605 214.415 ;
        RECT 51.105 212.415 52.105 213.415 ;
        RECT 53.605 212.415 54.605 213.415 ;
        RECT 51.105 211.415 54.605 212.415 ;
        RECT 55.605 213.415 59.105 214.415 ;
        RECT 60.105 213.415 63.605 214.415 ;
        RECT 46.605 209.415 50.105 210.415 ;
        RECT 51.105 209.415 52.105 211.415 ;
        RECT 55.605 210.415 56.605 213.415 ;
        RECT 60.105 212.415 61.105 213.415 ;
        RECT 62.605 212.415 63.605 213.415 ;
        RECT 60.105 211.415 63.605 212.415 ;
        RECT 64.605 213.415 68.105 214.415 ;
        RECT 64.605 212.415 65.605 213.415 ;
        RECT 64.605 211.415 68.105 212.415 ;
        RECT 70.105 211.415 72.605 212.415 ;
        RECT 55.605 209.415 59.105 210.415 ;
        RECT 60.105 209.415 61.105 211.415 ;
        RECT 62.605 209.415 63.605 211.415 ;
        RECT 67.105 210.415 68.105 211.415 ;
        RECT 64.605 209.415 68.105 210.415 ;
        RECT 73.605 209.415 74.605 214.415 ;
        RECT 75.605 209.415 76.605 214.415 ;
        RECT 77.605 213.415 81.605 214.415 ;
        RECT 82.605 213.415 86.605 214.415 ;
        RECT 87.605 213.915 88.605 214.415 ;
        RECT 79.105 209.415 80.105 213.415 ;
        RECT 82.605 210.415 83.605 213.415 ;
        RECT 87.605 212.915 89.605 213.915 ;
        RECT 84.605 211.415 86.605 212.415 ;
        RECT 85.605 210.415 86.605 211.415 ;
        RECT 82.605 209.415 86.605 210.415 ;
        RECT 87.605 209.415 88.605 212.915 ;
        RECT 89.105 212.415 90.105 212.915 ;
        RECT 89.605 211.915 90.605 212.415 ;
        RECT 90.105 211.415 91.105 211.915 ;
        RECT 91.605 211.415 92.605 214.415 ;
        RECT 90.605 210.915 92.605 211.415 ;
        RECT 91.105 210.415 92.605 210.915 ;
        RECT 91.605 209.415 92.605 210.415 ;
        RECT 42.730 203.750 43.230 204.250 ;
        RECT 42.730 203.250 43.730 203.750 ;
        RECT 42.730 202.750 44.230 203.250 ;
        RECT 42.730 200.750 43.230 202.750 ;
        RECT 43.730 202.250 44.730 202.750 ;
        RECT 45.230 202.250 45.730 204.250 ;
        RECT 44.230 201.750 45.730 202.250 ;
        RECT 44.730 201.250 45.730 201.750 ;
        RECT 45.230 200.750 45.730 201.250 ;
        RECT 46.230 200.750 46.730 204.250 ;
        RECT 47.230 203.750 49.730 204.250 ;
        RECT 48.230 200.750 48.730 203.750 ;
        RECT 50.230 202.750 50.730 204.250 ;
        RECT 52.230 202.750 52.730 204.250 ;
        RECT 50.230 202.250 52.730 202.750 ;
        RECT 50.230 200.750 50.730 202.250 ;
        RECT 52.230 200.750 52.730 202.250 ;
        RECT 53.230 200.750 53.730 204.250 ;
        RECT 54.230 203.750 54.730 204.250 ;
        RECT 54.230 203.250 55.230 203.750 ;
        RECT 54.230 202.750 55.730 203.250 ;
        RECT 54.230 200.750 54.730 202.750 ;
        RECT 55.230 202.250 56.230 202.750 ;
        RECT 56.730 202.250 57.230 204.250 ;
        RECT 55.730 201.750 57.230 202.250 ;
        RECT 56.230 201.250 57.230 201.750 ;
        RECT 56.730 200.750 57.230 201.250 ;
        RECT 58.230 203.750 60.230 204.250 ;
        RECT 58.230 202.750 58.730 203.750 ;
        RECT 59.730 202.750 60.230 203.750 ;
        RECT 58.230 202.250 60.230 202.750 ;
        RECT 62.730 202.750 63.230 204.250 ;
        RECT 64.730 203.750 65.230 204.250 ;
        RECT 64.230 203.250 65.230 203.750 ;
        RECT 65.730 203.750 67.730 204.250 ;
        RECT 63.730 202.750 64.730 203.250 ;
        RECT 65.730 202.750 66.230 203.750 ;
        RECT 67.230 202.750 67.730 203.750 ;
        RECT 62.730 202.250 64.230 202.750 ;
        RECT 65.730 202.250 67.730 202.750 ;
        RECT 58.230 200.750 58.730 202.250 ;
        RECT 62.730 200.750 63.230 202.250 ;
        RECT 63.730 201.750 64.730 202.250 ;
        RECT 64.230 201.250 65.230 201.750 ;
        RECT 64.730 200.750 65.230 201.250 ;
        RECT 65.730 200.750 66.230 202.250 ;
        RECT 67.230 200.750 67.730 202.250 ;
        RECT 68.230 203.750 70.230 204.250 ;
        RECT 70.730 203.750 73.230 204.250 ;
        RECT 68.230 202.750 68.730 203.750 ;
        RECT 69.730 202.750 70.230 203.750 ;
        RECT 68.230 202.250 70.230 202.750 ;
        RECT 68.230 200.750 68.730 202.250 ;
        RECT 69.230 201.750 69.730 202.250 ;
        RECT 69.230 201.250 70.230 201.750 ;
        RECT 69.730 200.750 70.230 201.250 ;
        RECT 71.730 200.750 72.230 203.750 ;
        RECT 73.730 200.750 74.230 204.250 ;
        RECT 74.730 202.750 75.230 204.250 ;
        RECT 76.730 203.750 77.230 204.250 ;
        RECT 76.230 203.250 77.230 203.750 ;
        RECT 77.730 203.750 79.730 204.250 ;
        RECT 75.730 202.750 76.730 203.250 ;
        RECT 77.730 202.750 78.230 203.750 ;
        RECT 79.230 202.750 79.730 203.750 ;
        RECT 74.730 202.250 76.230 202.750 ;
        RECT 77.730 202.250 79.730 202.750 ;
        RECT 80.230 202.750 80.730 204.250 ;
        RECT 81.730 202.750 82.230 204.250 ;
        RECT 80.230 202.250 82.230 202.750 ;
        RECT 84.730 203.750 85.730 204.250 ;
        RECT 87.230 203.750 88.230 204.250 ;
        RECT 84.730 203.250 86.230 203.750 ;
        RECT 86.730 203.250 88.230 203.750 ;
        RECT 74.730 200.750 75.230 202.250 ;
        RECT 75.730 201.750 76.730 202.250 ;
        RECT 76.230 201.250 77.230 201.750 ;
        RECT 76.730 200.750 77.230 201.250 ;
        RECT 77.730 200.750 78.230 202.250 ;
        RECT 79.230 200.750 79.730 202.250 ;
        RECT 80.980 200.750 81.480 202.250 ;
        RECT 84.730 200.750 85.230 203.250 ;
        RECT 85.730 202.750 88.230 203.250 ;
        RECT 86.230 202.250 86.730 202.750 ;
        RECT 87.730 200.750 88.230 202.750 ;
        RECT 88.730 203.750 90.730 204.250 ;
        RECT 88.730 202.750 89.230 203.750 ;
        RECT 90.230 202.750 90.730 203.750 ;
        RECT 88.730 202.250 90.730 202.750 ;
        RECT 88.730 200.750 89.230 202.250 ;
        RECT 90.230 200.750 90.730 202.250 ;
        RECT 91.230 203.750 93.230 204.250 ;
        RECT 91.230 201.250 91.730 203.750 ;
        RECT 92.730 203.250 93.730 203.750 ;
        RECT 93.230 201.750 93.730 203.250 ;
        RECT 92.730 201.250 93.730 201.750 ;
        RECT 94.230 202.750 94.730 204.250 ;
        RECT 95.730 202.750 96.230 204.250 ;
        RECT 94.230 202.250 96.230 202.750 ;
        RECT 91.230 200.750 93.230 201.250 ;
        RECT 94.230 200.750 94.730 202.250 ;
        RECT 95.730 200.750 96.230 202.250 ;
        RECT 96.730 203.750 98.730 204.250 ;
        RECT 96.730 202.750 97.230 203.750 ;
        RECT 98.230 202.750 98.730 203.750 ;
        RECT 96.730 202.250 98.730 202.750 ;
        RECT 96.730 200.750 97.230 202.250 ;
        RECT 98.230 200.750 98.730 202.250 ;
        RECT 99.230 202.250 99.730 204.250 ;
        RECT 101.730 202.250 102.230 204.250 ;
        RECT 99.230 201.750 100.230 202.250 ;
        RECT 101.230 201.750 102.230 202.250 ;
        RECT 103.230 203.750 105.730 204.250 ;
        RECT 103.230 202.750 103.730 203.750 ;
        RECT 104.730 202.750 105.730 203.750 ;
        RECT 103.230 202.250 105.730 202.750 ;
        RECT 99.730 201.250 101.730 201.750 ;
        RECT 100.230 200.750 101.230 201.250 ;
        RECT 103.230 200.750 103.730 202.250 ;
        RECT 114.390 192.310 114.690 224.760 ;
        RECT 42.830 191.700 114.690 192.310 ;
        RECT 42.830 191.650 114.680 191.700 ;
        RECT 42.830 191.640 45.470 191.650 ;
        RECT 117.150 189.360 117.450 224.760 ;
        RECT 37.390 188.790 117.450 189.360 ;
        RECT 9.200 166.970 26.930 167.390 ;
        RECT 37.400 165.490 37.980 188.790 ;
        RECT 36.780 165.180 106.430 165.190 ;
        RECT 116.780 165.180 118.940 168.290 ;
        RECT 36.780 165.170 118.940 165.180 ;
        RECT 36.780 164.610 118.910 165.170 ;
        RECT 36.640 61.500 38.230 62.680 ;
        RECT 39.570 4.920 40.470 164.610 ;
        RECT 45.040 158.410 45.500 158.420 ;
        RECT 45.040 8.000 45.830 158.410 ;
        RECT 82.170 156.920 93.470 156.940 ;
        RECT 81.630 155.250 93.470 156.920 ;
        RECT 81.640 154.620 82.150 155.250 ;
        RECT 76.105 153.625 76.625 154.620 ;
        RECT 72.435 151.010 80.295 153.625 ;
        RECT 49.920 148.920 80.295 151.010 ;
        RECT 72.435 145.765 80.295 148.920 ;
        RECT 76.105 143.775 76.625 145.765 ;
        RECT 72.435 135.915 80.295 143.775 ;
        RECT 76.105 133.925 76.625 135.915 ;
        RECT 72.435 126.065 80.295 133.925 ;
        RECT 76.105 124.075 76.625 126.065 ;
        RECT 72.435 116.215 80.295 124.075 ;
        RECT 76.105 115.480 76.625 116.215 ;
        RECT 76.100 114.300 76.630 115.480 ;
        RECT 81.630 115.220 82.150 154.620 ;
        RECT 87.415 153.625 87.935 154.620 ;
        RECT 92.940 154.020 93.470 155.250 ;
        RECT 83.745 145.765 91.605 153.625 ;
        RECT 87.415 143.775 87.935 145.765 ;
        RECT 83.745 135.915 91.605 143.775 ;
        RECT 87.415 133.925 87.935 135.915 ;
        RECT 83.745 126.065 91.605 133.925 ;
        RECT 87.415 124.075 87.935 126.065 ;
        RECT 83.745 116.215 91.605 124.075 ;
        RECT 87.415 115.700 87.935 116.215 ;
        RECT 87.410 114.300 87.940 115.700 ;
        RECT 92.940 115.220 93.460 154.020 ;
        RECT 76.100 113.830 87.940 114.300 ;
        RECT 52.910 99.920 53.430 99.940 ;
        RECT 119.910 99.920 120.210 224.760 ;
        RECT 52.910 99.420 120.210 99.920 ;
        RECT 122.670 98.130 122.970 224.760 ;
        RECT 47.480 97.610 122.970 98.130 ;
        RECT 47.480 91.020 47.980 97.610 ;
        RECT 136.170 95.680 137.070 96.900 ;
        RECT 128.570 95.190 137.070 95.680 ;
        RECT 47.480 73.630 48.010 91.020 ;
        RECT 52.920 76.010 53.410 76.560 ;
        RECT 46.840 73.300 116.490 73.310 ;
        RECT 126.840 73.300 129.000 76.410 ;
        RECT 46.840 73.290 129.000 73.300 ;
        RECT 46.840 72.730 128.970 73.290 ;
        RECT 54.310 10.270 54.830 69.120 ;
        RECT 97.530 65.060 98.430 72.730 ;
        RECT 92.230 65.040 103.530 65.060 ;
        RECT 91.690 63.370 103.530 65.040 ;
        RECT 91.700 62.740 92.210 63.370 ;
        RECT 97.530 62.740 98.430 63.370 ;
        RECT 86.165 61.745 86.685 62.740 ;
        RECT 82.495 59.130 90.355 61.745 ;
        RECT 59.980 57.040 90.355 59.130 ;
        RECT 82.495 53.885 90.355 57.040 ;
        RECT 86.165 51.895 86.685 53.885 ;
        RECT 82.495 44.035 90.355 51.895 ;
        RECT 86.165 42.045 86.685 44.035 ;
        RECT 82.495 34.185 90.355 42.045 ;
        RECT 86.165 32.195 86.685 34.185 ;
        RECT 82.495 24.335 90.355 32.195 ;
        RECT 86.165 23.600 86.685 24.335 ;
        RECT 86.160 22.420 86.690 23.600 ;
        RECT 91.690 23.340 92.210 62.740 ;
        RECT 97.475 61.745 98.430 62.740 ;
        RECT 103.000 62.140 103.530 63.370 ;
        RECT 93.805 53.885 101.665 61.745 ;
        RECT 97.475 51.895 98.430 53.885 ;
        RECT 93.805 44.035 101.665 51.895 ;
        RECT 97.475 42.045 98.430 44.035 ;
        RECT 93.805 34.185 101.665 42.045 ;
        RECT 97.475 32.195 98.430 34.185 ;
        RECT 93.805 24.335 101.665 32.195 ;
        RECT 97.475 23.820 98.430 24.335 ;
        RECT 97.470 22.420 98.430 23.820 ;
        RECT 103.000 23.340 103.520 62.140 ;
        RECT 86.160 21.950 98.430 22.420 ;
        RECT 54.300 9.150 98.430 10.270 ;
        RECT 54.300 9.140 56.070 9.150 ;
        RECT 77.840 8.000 79.110 8.010 ;
        RECT 45.040 7.990 56.100 8.000 ;
        RECT 60.800 7.990 79.110 8.000 ;
        RECT 45.040 7.100 79.110 7.990 ;
        RECT 45.950 4.920 59.790 4.930 ;
        RECT 39.560 4.120 59.790 4.920 ;
        RECT 45.950 4.100 59.790 4.120 ;
        RECT 58.890 1.000 59.790 4.100 ;
        RECT 78.210 1.000 79.110 7.100 ;
        RECT 97.530 1.000 98.430 9.150 ;
        RECT 116.850 1.000 117.750 72.730 ;
        RECT 136.170 1.000 137.070 95.190 ;
  END
END tt_um_LPCAS_TP1
END LIBRARY

