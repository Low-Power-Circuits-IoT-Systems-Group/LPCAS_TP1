magic
tech sky130A
magscale 1 2
timestamp 1741700111
<< locali >>
rect -19 -17 19 17
<< viali >>
rect -53 -17 -19 17
rect 19 -17 53 17
<< metal1 >>
rect -68 17 68 23
rect -68 -17 -53 17
rect -19 -17 19 17
rect 53 -17 68 17
rect -68 -23 68 -17
<< end >>
